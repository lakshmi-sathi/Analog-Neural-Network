magic
tech sky130A
magscale 1 2
timestamp 1627812032
<< pwell >>
rect -360 -648 360 648
<< psubdiff >>
rect -324 578 -228 612
rect 228 578 324 612
rect -324 516 -290 578
rect 290 516 324 578
rect -324 -578 -290 -516
rect 290 -578 324 -516
rect -324 -612 -228 -578
rect 228 -612 324 -578
<< psubdiffcont >>
rect -228 578 228 612
rect -324 -516 -290 516
rect 290 -516 324 516
rect -228 -612 228 -578
<< xpolycontact >>
rect -194 50 -124 482
rect -194 -482 -124 -50
rect 124 50 194 482
rect 124 -482 194 -50
<< ppolyres >>
rect -194 -50 -124 50
rect 124 -50 194 50
<< locali >>
rect -324 578 -228 612
rect 228 578 324 612
rect -324 516 -290 578
rect 290 516 324 578
rect -324 -578 -290 -516
rect 290 -578 324 -516
rect -324 -612 -228 -578
rect 228 -612 324 -578
<< viali >>
rect -178 67 -140 464
rect 140 67 178 464
rect -178 -464 -140 -67
rect 140 -464 178 -67
<< metal1 >>
rect -184 464 -134 476
rect -184 67 -178 464
rect -140 67 -134 464
rect -184 55 -134 67
rect 134 464 184 476
rect 134 67 140 464
rect 178 67 184 464
rect 134 55 184 67
rect -184 -67 -134 -55
rect -184 -464 -178 -67
rect -140 -464 -134 -67
rect -184 -476 -134 -464
rect 134 -67 184 -55
rect 134 -464 140 -67
rect 178 -464 184 -67
rect 134 -476 184 -464
<< res0p35 >>
rect -196 -52 -122 52
rect 122 -52 196 52
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string FIXED_BBOX -307 -595 307 595
string parameters w 0.350 l 0.50 m 1 nx 2 wmin 0.350 lmin 0.50 rho 319.8 val 566.502 dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
