magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_p >>
rect -845 641 -787 647
rect -653 641 -595 647
rect -461 641 -403 647
rect -269 641 -211 647
rect -77 641 -19 647
rect 115 641 173 647
rect 307 641 365 647
rect 499 641 557 647
rect 691 641 749 647
rect -845 607 -833 641
rect -653 607 -641 641
rect -461 607 -449 641
rect -269 607 -257 641
rect -77 607 -65 641
rect 115 607 127 641
rect 307 607 319 641
rect 499 607 511 641
rect 691 607 703 641
rect -845 601 -787 607
rect -653 601 -595 607
rect -461 601 -403 607
rect -269 601 -211 607
rect -77 601 -19 607
rect 115 601 173 607
rect 307 601 365 607
rect 499 601 557 607
rect 691 601 749 607
rect -749 71 -691 77
rect -557 71 -499 77
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect 595 71 653 77
rect 787 71 845 77
rect -749 37 -737 71
rect -557 37 -545 71
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect 595 37 607 71
rect 787 37 799 71
rect -749 31 -691 37
rect -557 31 -499 37
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect 595 31 653 37
rect 787 31 845 37
rect -749 -37 -691 -31
rect -557 -37 -499 -31
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect 595 -37 653 -31
rect 787 -37 845 -31
rect -749 -71 -737 -37
rect -557 -71 -545 -37
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect 595 -71 607 -37
rect 787 -71 799 -37
rect -749 -77 -691 -71
rect -557 -77 -499 -71
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect 595 -77 653 -71
rect 787 -77 845 -71
rect -845 -607 -787 -601
rect -653 -607 -595 -601
rect -461 -607 -403 -601
rect -269 -607 -211 -601
rect -77 -607 -19 -601
rect 115 -607 173 -601
rect 307 -607 365 -601
rect 499 -607 557 -601
rect 691 -607 749 -601
rect -845 -641 -833 -607
rect -653 -641 -641 -607
rect -461 -641 -449 -607
rect -269 -641 -257 -607
rect -77 -641 -65 -607
rect 115 -641 127 -607
rect 307 -641 319 -607
rect 499 -641 511 -607
rect 691 -641 703 -607
rect -845 -647 -787 -641
rect -653 -647 -595 -641
rect -461 -647 -403 -641
rect -269 -647 -211 -641
rect -77 -647 -19 -641
rect 115 -647 173 -641
rect 307 -647 365 -641
rect 499 -647 557 -641
rect 691 -647 749 -641
<< nwell >>
rect -1031 -779 1031 779
<< pmos >>
rect -831 118 -801 560
rect -735 118 -705 560
rect -639 118 -609 560
rect -543 118 -513 560
rect -447 118 -417 560
rect -351 118 -321 560
rect -255 118 -225 560
rect -159 118 -129 560
rect -63 118 -33 560
rect 33 118 63 560
rect 129 118 159 560
rect 225 118 255 560
rect 321 118 351 560
rect 417 118 447 560
rect 513 118 543 560
rect 609 118 639 560
rect 705 118 735 560
rect 801 118 831 560
rect -831 -560 -801 -118
rect -735 -560 -705 -118
rect -639 -560 -609 -118
rect -543 -560 -513 -118
rect -447 -560 -417 -118
rect -351 -560 -321 -118
rect -255 -560 -225 -118
rect -159 -560 -129 -118
rect -63 -560 -33 -118
rect 33 -560 63 -118
rect 129 -560 159 -118
rect 225 -560 255 -118
rect 321 -560 351 -118
rect 417 -560 447 -118
rect 513 -560 543 -118
rect 609 -560 639 -118
rect 705 -560 735 -118
rect 801 -560 831 -118
<< pdiff >>
rect -893 526 -831 560
rect -893 492 -881 526
rect -847 492 -831 526
rect -893 458 -831 492
rect -893 424 -881 458
rect -847 424 -831 458
rect -893 390 -831 424
rect -893 356 -881 390
rect -847 356 -831 390
rect -893 322 -831 356
rect -893 288 -881 322
rect -847 288 -831 322
rect -893 254 -831 288
rect -893 220 -881 254
rect -847 220 -831 254
rect -893 186 -831 220
rect -893 152 -881 186
rect -847 152 -831 186
rect -893 118 -831 152
rect -801 526 -735 560
rect -801 492 -785 526
rect -751 492 -735 526
rect -801 458 -735 492
rect -801 424 -785 458
rect -751 424 -735 458
rect -801 390 -735 424
rect -801 356 -785 390
rect -751 356 -735 390
rect -801 322 -735 356
rect -801 288 -785 322
rect -751 288 -735 322
rect -801 254 -735 288
rect -801 220 -785 254
rect -751 220 -735 254
rect -801 186 -735 220
rect -801 152 -785 186
rect -751 152 -735 186
rect -801 118 -735 152
rect -705 526 -639 560
rect -705 492 -689 526
rect -655 492 -639 526
rect -705 458 -639 492
rect -705 424 -689 458
rect -655 424 -639 458
rect -705 390 -639 424
rect -705 356 -689 390
rect -655 356 -639 390
rect -705 322 -639 356
rect -705 288 -689 322
rect -655 288 -639 322
rect -705 254 -639 288
rect -705 220 -689 254
rect -655 220 -639 254
rect -705 186 -639 220
rect -705 152 -689 186
rect -655 152 -639 186
rect -705 118 -639 152
rect -609 526 -543 560
rect -609 492 -593 526
rect -559 492 -543 526
rect -609 458 -543 492
rect -609 424 -593 458
rect -559 424 -543 458
rect -609 390 -543 424
rect -609 356 -593 390
rect -559 356 -543 390
rect -609 322 -543 356
rect -609 288 -593 322
rect -559 288 -543 322
rect -609 254 -543 288
rect -609 220 -593 254
rect -559 220 -543 254
rect -609 186 -543 220
rect -609 152 -593 186
rect -559 152 -543 186
rect -609 118 -543 152
rect -513 526 -447 560
rect -513 492 -497 526
rect -463 492 -447 526
rect -513 458 -447 492
rect -513 424 -497 458
rect -463 424 -447 458
rect -513 390 -447 424
rect -513 356 -497 390
rect -463 356 -447 390
rect -513 322 -447 356
rect -513 288 -497 322
rect -463 288 -447 322
rect -513 254 -447 288
rect -513 220 -497 254
rect -463 220 -447 254
rect -513 186 -447 220
rect -513 152 -497 186
rect -463 152 -447 186
rect -513 118 -447 152
rect -417 526 -351 560
rect -417 492 -401 526
rect -367 492 -351 526
rect -417 458 -351 492
rect -417 424 -401 458
rect -367 424 -351 458
rect -417 390 -351 424
rect -417 356 -401 390
rect -367 356 -351 390
rect -417 322 -351 356
rect -417 288 -401 322
rect -367 288 -351 322
rect -417 254 -351 288
rect -417 220 -401 254
rect -367 220 -351 254
rect -417 186 -351 220
rect -417 152 -401 186
rect -367 152 -351 186
rect -417 118 -351 152
rect -321 526 -255 560
rect -321 492 -305 526
rect -271 492 -255 526
rect -321 458 -255 492
rect -321 424 -305 458
rect -271 424 -255 458
rect -321 390 -255 424
rect -321 356 -305 390
rect -271 356 -255 390
rect -321 322 -255 356
rect -321 288 -305 322
rect -271 288 -255 322
rect -321 254 -255 288
rect -321 220 -305 254
rect -271 220 -255 254
rect -321 186 -255 220
rect -321 152 -305 186
rect -271 152 -255 186
rect -321 118 -255 152
rect -225 526 -159 560
rect -225 492 -209 526
rect -175 492 -159 526
rect -225 458 -159 492
rect -225 424 -209 458
rect -175 424 -159 458
rect -225 390 -159 424
rect -225 356 -209 390
rect -175 356 -159 390
rect -225 322 -159 356
rect -225 288 -209 322
rect -175 288 -159 322
rect -225 254 -159 288
rect -225 220 -209 254
rect -175 220 -159 254
rect -225 186 -159 220
rect -225 152 -209 186
rect -175 152 -159 186
rect -225 118 -159 152
rect -129 526 -63 560
rect -129 492 -113 526
rect -79 492 -63 526
rect -129 458 -63 492
rect -129 424 -113 458
rect -79 424 -63 458
rect -129 390 -63 424
rect -129 356 -113 390
rect -79 356 -63 390
rect -129 322 -63 356
rect -129 288 -113 322
rect -79 288 -63 322
rect -129 254 -63 288
rect -129 220 -113 254
rect -79 220 -63 254
rect -129 186 -63 220
rect -129 152 -113 186
rect -79 152 -63 186
rect -129 118 -63 152
rect -33 526 33 560
rect -33 492 -17 526
rect 17 492 33 526
rect -33 458 33 492
rect -33 424 -17 458
rect 17 424 33 458
rect -33 390 33 424
rect -33 356 -17 390
rect 17 356 33 390
rect -33 322 33 356
rect -33 288 -17 322
rect 17 288 33 322
rect -33 254 33 288
rect -33 220 -17 254
rect 17 220 33 254
rect -33 186 33 220
rect -33 152 -17 186
rect 17 152 33 186
rect -33 118 33 152
rect 63 526 129 560
rect 63 492 79 526
rect 113 492 129 526
rect 63 458 129 492
rect 63 424 79 458
rect 113 424 129 458
rect 63 390 129 424
rect 63 356 79 390
rect 113 356 129 390
rect 63 322 129 356
rect 63 288 79 322
rect 113 288 129 322
rect 63 254 129 288
rect 63 220 79 254
rect 113 220 129 254
rect 63 186 129 220
rect 63 152 79 186
rect 113 152 129 186
rect 63 118 129 152
rect 159 526 225 560
rect 159 492 175 526
rect 209 492 225 526
rect 159 458 225 492
rect 159 424 175 458
rect 209 424 225 458
rect 159 390 225 424
rect 159 356 175 390
rect 209 356 225 390
rect 159 322 225 356
rect 159 288 175 322
rect 209 288 225 322
rect 159 254 225 288
rect 159 220 175 254
rect 209 220 225 254
rect 159 186 225 220
rect 159 152 175 186
rect 209 152 225 186
rect 159 118 225 152
rect 255 526 321 560
rect 255 492 271 526
rect 305 492 321 526
rect 255 458 321 492
rect 255 424 271 458
rect 305 424 321 458
rect 255 390 321 424
rect 255 356 271 390
rect 305 356 321 390
rect 255 322 321 356
rect 255 288 271 322
rect 305 288 321 322
rect 255 254 321 288
rect 255 220 271 254
rect 305 220 321 254
rect 255 186 321 220
rect 255 152 271 186
rect 305 152 321 186
rect 255 118 321 152
rect 351 526 417 560
rect 351 492 367 526
rect 401 492 417 526
rect 351 458 417 492
rect 351 424 367 458
rect 401 424 417 458
rect 351 390 417 424
rect 351 356 367 390
rect 401 356 417 390
rect 351 322 417 356
rect 351 288 367 322
rect 401 288 417 322
rect 351 254 417 288
rect 351 220 367 254
rect 401 220 417 254
rect 351 186 417 220
rect 351 152 367 186
rect 401 152 417 186
rect 351 118 417 152
rect 447 526 513 560
rect 447 492 463 526
rect 497 492 513 526
rect 447 458 513 492
rect 447 424 463 458
rect 497 424 513 458
rect 447 390 513 424
rect 447 356 463 390
rect 497 356 513 390
rect 447 322 513 356
rect 447 288 463 322
rect 497 288 513 322
rect 447 254 513 288
rect 447 220 463 254
rect 497 220 513 254
rect 447 186 513 220
rect 447 152 463 186
rect 497 152 513 186
rect 447 118 513 152
rect 543 526 609 560
rect 543 492 559 526
rect 593 492 609 526
rect 543 458 609 492
rect 543 424 559 458
rect 593 424 609 458
rect 543 390 609 424
rect 543 356 559 390
rect 593 356 609 390
rect 543 322 609 356
rect 543 288 559 322
rect 593 288 609 322
rect 543 254 609 288
rect 543 220 559 254
rect 593 220 609 254
rect 543 186 609 220
rect 543 152 559 186
rect 593 152 609 186
rect 543 118 609 152
rect 639 526 705 560
rect 639 492 655 526
rect 689 492 705 526
rect 639 458 705 492
rect 639 424 655 458
rect 689 424 705 458
rect 639 390 705 424
rect 639 356 655 390
rect 689 356 705 390
rect 639 322 705 356
rect 639 288 655 322
rect 689 288 705 322
rect 639 254 705 288
rect 639 220 655 254
rect 689 220 705 254
rect 639 186 705 220
rect 639 152 655 186
rect 689 152 705 186
rect 639 118 705 152
rect 735 526 801 560
rect 735 492 751 526
rect 785 492 801 526
rect 735 458 801 492
rect 735 424 751 458
rect 785 424 801 458
rect 735 390 801 424
rect 735 356 751 390
rect 785 356 801 390
rect 735 322 801 356
rect 735 288 751 322
rect 785 288 801 322
rect 735 254 801 288
rect 735 220 751 254
rect 785 220 801 254
rect 735 186 801 220
rect 735 152 751 186
rect 785 152 801 186
rect 735 118 801 152
rect 831 526 893 560
rect 831 492 847 526
rect 881 492 893 526
rect 831 458 893 492
rect 831 424 847 458
rect 881 424 893 458
rect 831 390 893 424
rect 831 356 847 390
rect 881 356 893 390
rect 831 322 893 356
rect 831 288 847 322
rect 881 288 893 322
rect 831 254 893 288
rect 831 220 847 254
rect 881 220 893 254
rect 831 186 893 220
rect 831 152 847 186
rect 881 152 893 186
rect 831 118 893 152
rect -893 -152 -831 -118
rect -893 -186 -881 -152
rect -847 -186 -831 -152
rect -893 -220 -831 -186
rect -893 -254 -881 -220
rect -847 -254 -831 -220
rect -893 -288 -831 -254
rect -893 -322 -881 -288
rect -847 -322 -831 -288
rect -893 -356 -831 -322
rect -893 -390 -881 -356
rect -847 -390 -831 -356
rect -893 -424 -831 -390
rect -893 -458 -881 -424
rect -847 -458 -831 -424
rect -893 -492 -831 -458
rect -893 -526 -881 -492
rect -847 -526 -831 -492
rect -893 -560 -831 -526
rect -801 -152 -735 -118
rect -801 -186 -785 -152
rect -751 -186 -735 -152
rect -801 -220 -735 -186
rect -801 -254 -785 -220
rect -751 -254 -735 -220
rect -801 -288 -735 -254
rect -801 -322 -785 -288
rect -751 -322 -735 -288
rect -801 -356 -735 -322
rect -801 -390 -785 -356
rect -751 -390 -735 -356
rect -801 -424 -735 -390
rect -801 -458 -785 -424
rect -751 -458 -735 -424
rect -801 -492 -735 -458
rect -801 -526 -785 -492
rect -751 -526 -735 -492
rect -801 -560 -735 -526
rect -705 -152 -639 -118
rect -705 -186 -689 -152
rect -655 -186 -639 -152
rect -705 -220 -639 -186
rect -705 -254 -689 -220
rect -655 -254 -639 -220
rect -705 -288 -639 -254
rect -705 -322 -689 -288
rect -655 -322 -639 -288
rect -705 -356 -639 -322
rect -705 -390 -689 -356
rect -655 -390 -639 -356
rect -705 -424 -639 -390
rect -705 -458 -689 -424
rect -655 -458 -639 -424
rect -705 -492 -639 -458
rect -705 -526 -689 -492
rect -655 -526 -639 -492
rect -705 -560 -639 -526
rect -609 -152 -543 -118
rect -609 -186 -593 -152
rect -559 -186 -543 -152
rect -609 -220 -543 -186
rect -609 -254 -593 -220
rect -559 -254 -543 -220
rect -609 -288 -543 -254
rect -609 -322 -593 -288
rect -559 -322 -543 -288
rect -609 -356 -543 -322
rect -609 -390 -593 -356
rect -559 -390 -543 -356
rect -609 -424 -543 -390
rect -609 -458 -593 -424
rect -559 -458 -543 -424
rect -609 -492 -543 -458
rect -609 -526 -593 -492
rect -559 -526 -543 -492
rect -609 -560 -543 -526
rect -513 -152 -447 -118
rect -513 -186 -497 -152
rect -463 -186 -447 -152
rect -513 -220 -447 -186
rect -513 -254 -497 -220
rect -463 -254 -447 -220
rect -513 -288 -447 -254
rect -513 -322 -497 -288
rect -463 -322 -447 -288
rect -513 -356 -447 -322
rect -513 -390 -497 -356
rect -463 -390 -447 -356
rect -513 -424 -447 -390
rect -513 -458 -497 -424
rect -463 -458 -447 -424
rect -513 -492 -447 -458
rect -513 -526 -497 -492
rect -463 -526 -447 -492
rect -513 -560 -447 -526
rect -417 -152 -351 -118
rect -417 -186 -401 -152
rect -367 -186 -351 -152
rect -417 -220 -351 -186
rect -417 -254 -401 -220
rect -367 -254 -351 -220
rect -417 -288 -351 -254
rect -417 -322 -401 -288
rect -367 -322 -351 -288
rect -417 -356 -351 -322
rect -417 -390 -401 -356
rect -367 -390 -351 -356
rect -417 -424 -351 -390
rect -417 -458 -401 -424
rect -367 -458 -351 -424
rect -417 -492 -351 -458
rect -417 -526 -401 -492
rect -367 -526 -351 -492
rect -417 -560 -351 -526
rect -321 -152 -255 -118
rect -321 -186 -305 -152
rect -271 -186 -255 -152
rect -321 -220 -255 -186
rect -321 -254 -305 -220
rect -271 -254 -255 -220
rect -321 -288 -255 -254
rect -321 -322 -305 -288
rect -271 -322 -255 -288
rect -321 -356 -255 -322
rect -321 -390 -305 -356
rect -271 -390 -255 -356
rect -321 -424 -255 -390
rect -321 -458 -305 -424
rect -271 -458 -255 -424
rect -321 -492 -255 -458
rect -321 -526 -305 -492
rect -271 -526 -255 -492
rect -321 -560 -255 -526
rect -225 -152 -159 -118
rect -225 -186 -209 -152
rect -175 -186 -159 -152
rect -225 -220 -159 -186
rect -225 -254 -209 -220
rect -175 -254 -159 -220
rect -225 -288 -159 -254
rect -225 -322 -209 -288
rect -175 -322 -159 -288
rect -225 -356 -159 -322
rect -225 -390 -209 -356
rect -175 -390 -159 -356
rect -225 -424 -159 -390
rect -225 -458 -209 -424
rect -175 -458 -159 -424
rect -225 -492 -159 -458
rect -225 -526 -209 -492
rect -175 -526 -159 -492
rect -225 -560 -159 -526
rect -129 -152 -63 -118
rect -129 -186 -113 -152
rect -79 -186 -63 -152
rect -129 -220 -63 -186
rect -129 -254 -113 -220
rect -79 -254 -63 -220
rect -129 -288 -63 -254
rect -129 -322 -113 -288
rect -79 -322 -63 -288
rect -129 -356 -63 -322
rect -129 -390 -113 -356
rect -79 -390 -63 -356
rect -129 -424 -63 -390
rect -129 -458 -113 -424
rect -79 -458 -63 -424
rect -129 -492 -63 -458
rect -129 -526 -113 -492
rect -79 -526 -63 -492
rect -129 -560 -63 -526
rect -33 -152 33 -118
rect -33 -186 -17 -152
rect 17 -186 33 -152
rect -33 -220 33 -186
rect -33 -254 -17 -220
rect 17 -254 33 -220
rect -33 -288 33 -254
rect -33 -322 -17 -288
rect 17 -322 33 -288
rect -33 -356 33 -322
rect -33 -390 -17 -356
rect 17 -390 33 -356
rect -33 -424 33 -390
rect -33 -458 -17 -424
rect 17 -458 33 -424
rect -33 -492 33 -458
rect -33 -526 -17 -492
rect 17 -526 33 -492
rect -33 -560 33 -526
rect 63 -152 129 -118
rect 63 -186 79 -152
rect 113 -186 129 -152
rect 63 -220 129 -186
rect 63 -254 79 -220
rect 113 -254 129 -220
rect 63 -288 129 -254
rect 63 -322 79 -288
rect 113 -322 129 -288
rect 63 -356 129 -322
rect 63 -390 79 -356
rect 113 -390 129 -356
rect 63 -424 129 -390
rect 63 -458 79 -424
rect 113 -458 129 -424
rect 63 -492 129 -458
rect 63 -526 79 -492
rect 113 -526 129 -492
rect 63 -560 129 -526
rect 159 -152 225 -118
rect 159 -186 175 -152
rect 209 -186 225 -152
rect 159 -220 225 -186
rect 159 -254 175 -220
rect 209 -254 225 -220
rect 159 -288 225 -254
rect 159 -322 175 -288
rect 209 -322 225 -288
rect 159 -356 225 -322
rect 159 -390 175 -356
rect 209 -390 225 -356
rect 159 -424 225 -390
rect 159 -458 175 -424
rect 209 -458 225 -424
rect 159 -492 225 -458
rect 159 -526 175 -492
rect 209 -526 225 -492
rect 159 -560 225 -526
rect 255 -152 321 -118
rect 255 -186 271 -152
rect 305 -186 321 -152
rect 255 -220 321 -186
rect 255 -254 271 -220
rect 305 -254 321 -220
rect 255 -288 321 -254
rect 255 -322 271 -288
rect 305 -322 321 -288
rect 255 -356 321 -322
rect 255 -390 271 -356
rect 305 -390 321 -356
rect 255 -424 321 -390
rect 255 -458 271 -424
rect 305 -458 321 -424
rect 255 -492 321 -458
rect 255 -526 271 -492
rect 305 -526 321 -492
rect 255 -560 321 -526
rect 351 -152 417 -118
rect 351 -186 367 -152
rect 401 -186 417 -152
rect 351 -220 417 -186
rect 351 -254 367 -220
rect 401 -254 417 -220
rect 351 -288 417 -254
rect 351 -322 367 -288
rect 401 -322 417 -288
rect 351 -356 417 -322
rect 351 -390 367 -356
rect 401 -390 417 -356
rect 351 -424 417 -390
rect 351 -458 367 -424
rect 401 -458 417 -424
rect 351 -492 417 -458
rect 351 -526 367 -492
rect 401 -526 417 -492
rect 351 -560 417 -526
rect 447 -152 513 -118
rect 447 -186 463 -152
rect 497 -186 513 -152
rect 447 -220 513 -186
rect 447 -254 463 -220
rect 497 -254 513 -220
rect 447 -288 513 -254
rect 447 -322 463 -288
rect 497 -322 513 -288
rect 447 -356 513 -322
rect 447 -390 463 -356
rect 497 -390 513 -356
rect 447 -424 513 -390
rect 447 -458 463 -424
rect 497 -458 513 -424
rect 447 -492 513 -458
rect 447 -526 463 -492
rect 497 -526 513 -492
rect 447 -560 513 -526
rect 543 -152 609 -118
rect 543 -186 559 -152
rect 593 -186 609 -152
rect 543 -220 609 -186
rect 543 -254 559 -220
rect 593 -254 609 -220
rect 543 -288 609 -254
rect 543 -322 559 -288
rect 593 -322 609 -288
rect 543 -356 609 -322
rect 543 -390 559 -356
rect 593 -390 609 -356
rect 543 -424 609 -390
rect 543 -458 559 -424
rect 593 -458 609 -424
rect 543 -492 609 -458
rect 543 -526 559 -492
rect 593 -526 609 -492
rect 543 -560 609 -526
rect 639 -152 705 -118
rect 639 -186 655 -152
rect 689 -186 705 -152
rect 639 -220 705 -186
rect 639 -254 655 -220
rect 689 -254 705 -220
rect 639 -288 705 -254
rect 639 -322 655 -288
rect 689 -322 705 -288
rect 639 -356 705 -322
rect 639 -390 655 -356
rect 689 -390 705 -356
rect 639 -424 705 -390
rect 639 -458 655 -424
rect 689 -458 705 -424
rect 639 -492 705 -458
rect 639 -526 655 -492
rect 689 -526 705 -492
rect 639 -560 705 -526
rect 735 -152 801 -118
rect 735 -186 751 -152
rect 785 -186 801 -152
rect 735 -220 801 -186
rect 735 -254 751 -220
rect 785 -254 801 -220
rect 735 -288 801 -254
rect 735 -322 751 -288
rect 785 -322 801 -288
rect 735 -356 801 -322
rect 735 -390 751 -356
rect 785 -390 801 -356
rect 735 -424 801 -390
rect 735 -458 751 -424
rect 785 -458 801 -424
rect 735 -492 801 -458
rect 735 -526 751 -492
rect 785 -526 801 -492
rect 735 -560 801 -526
rect 831 -152 893 -118
rect 831 -186 847 -152
rect 881 -186 893 -152
rect 831 -220 893 -186
rect 831 -254 847 -220
rect 881 -254 893 -220
rect 831 -288 893 -254
rect 831 -322 847 -288
rect 881 -322 893 -288
rect 831 -356 893 -322
rect 831 -390 847 -356
rect 881 -390 893 -356
rect 831 -424 893 -390
rect 831 -458 847 -424
rect 881 -458 893 -424
rect 831 -492 893 -458
rect 831 -526 847 -492
rect 881 -526 893 -492
rect 831 -560 893 -526
<< pdiffc >>
rect -881 492 -847 526
rect -881 424 -847 458
rect -881 356 -847 390
rect -881 288 -847 322
rect -881 220 -847 254
rect -881 152 -847 186
rect -785 492 -751 526
rect -785 424 -751 458
rect -785 356 -751 390
rect -785 288 -751 322
rect -785 220 -751 254
rect -785 152 -751 186
rect -689 492 -655 526
rect -689 424 -655 458
rect -689 356 -655 390
rect -689 288 -655 322
rect -689 220 -655 254
rect -689 152 -655 186
rect -593 492 -559 526
rect -593 424 -559 458
rect -593 356 -559 390
rect -593 288 -559 322
rect -593 220 -559 254
rect -593 152 -559 186
rect -497 492 -463 526
rect -497 424 -463 458
rect -497 356 -463 390
rect -497 288 -463 322
rect -497 220 -463 254
rect -497 152 -463 186
rect -401 492 -367 526
rect -401 424 -367 458
rect -401 356 -367 390
rect -401 288 -367 322
rect -401 220 -367 254
rect -401 152 -367 186
rect -305 492 -271 526
rect -305 424 -271 458
rect -305 356 -271 390
rect -305 288 -271 322
rect -305 220 -271 254
rect -305 152 -271 186
rect -209 492 -175 526
rect -209 424 -175 458
rect -209 356 -175 390
rect -209 288 -175 322
rect -209 220 -175 254
rect -209 152 -175 186
rect -113 492 -79 526
rect -113 424 -79 458
rect -113 356 -79 390
rect -113 288 -79 322
rect -113 220 -79 254
rect -113 152 -79 186
rect -17 492 17 526
rect -17 424 17 458
rect -17 356 17 390
rect -17 288 17 322
rect -17 220 17 254
rect -17 152 17 186
rect 79 492 113 526
rect 79 424 113 458
rect 79 356 113 390
rect 79 288 113 322
rect 79 220 113 254
rect 79 152 113 186
rect 175 492 209 526
rect 175 424 209 458
rect 175 356 209 390
rect 175 288 209 322
rect 175 220 209 254
rect 175 152 209 186
rect 271 492 305 526
rect 271 424 305 458
rect 271 356 305 390
rect 271 288 305 322
rect 271 220 305 254
rect 271 152 305 186
rect 367 492 401 526
rect 367 424 401 458
rect 367 356 401 390
rect 367 288 401 322
rect 367 220 401 254
rect 367 152 401 186
rect 463 492 497 526
rect 463 424 497 458
rect 463 356 497 390
rect 463 288 497 322
rect 463 220 497 254
rect 463 152 497 186
rect 559 492 593 526
rect 559 424 593 458
rect 559 356 593 390
rect 559 288 593 322
rect 559 220 593 254
rect 559 152 593 186
rect 655 492 689 526
rect 655 424 689 458
rect 655 356 689 390
rect 655 288 689 322
rect 655 220 689 254
rect 655 152 689 186
rect 751 492 785 526
rect 751 424 785 458
rect 751 356 785 390
rect 751 288 785 322
rect 751 220 785 254
rect 751 152 785 186
rect 847 492 881 526
rect 847 424 881 458
rect 847 356 881 390
rect 847 288 881 322
rect 847 220 881 254
rect 847 152 881 186
rect -881 -186 -847 -152
rect -881 -254 -847 -220
rect -881 -322 -847 -288
rect -881 -390 -847 -356
rect -881 -458 -847 -424
rect -881 -526 -847 -492
rect -785 -186 -751 -152
rect -785 -254 -751 -220
rect -785 -322 -751 -288
rect -785 -390 -751 -356
rect -785 -458 -751 -424
rect -785 -526 -751 -492
rect -689 -186 -655 -152
rect -689 -254 -655 -220
rect -689 -322 -655 -288
rect -689 -390 -655 -356
rect -689 -458 -655 -424
rect -689 -526 -655 -492
rect -593 -186 -559 -152
rect -593 -254 -559 -220
rect -593 -322 -559 -288
rect -593 -390 -559 -356
rect -593 -458 -559 -424
rect -593 -526 -559 -492
rect -497 -186 -463 -152
rect -497 -254 -463 -220
rect -497 -322 -463 -288
rect -497 -390 -463 -356
rect -497 -458 -463 -424
rect -497 -526 -463 -492
rect -401 -186 -367 -152
rect -401 -254 -367 -220
rect -401 -322 -367 -288
rect -401 -390 -367 -356
rect -401 -458 -367 -424
rect -401 -526 -367 -492
rect -305 -186 -271 -152
rect -305 -254 -271 -220
rect -305 -322 -271 -288
rect -305 -390 -271 -356
rect -305 -458 -271 -424
rect -305 -526 -271 -492
rect -209 -186 -175 -152
rect -209 -254 -175 -220
rect -209 -322 -175 -288
rect -209 -390 -175 -356
rect -209 -458 -175 -424
rect -209 -526 -175 -492
rect -113 -186 -79 -152
rect -113 -254 -79 -220
rect -113 -322 -79 -288
rect -113 -390 -79 -356
rect -113 -458 -79 -424
rect -113 -526 -79 -492
rect -17 -186 17 -152
rect -17 -254 17 -220
rect -17 -322 17 -288
rect -17 -390 17 -356
rect -17 -458 17 -424
rect -17 -526 17 -492
rect 79 -186 113 -152
rect 79 -254 113 -220
rect 79 -322 113 -288
rect 79 -390 113 -356
rect 79 -458 113 -424
rect 79 -526 113 -492
rect 175 -186 209 -152
rect 175 -254 209 -220
rect 175 -322 209 -288
rect 175 -390 209 -356
rect 175 -458 209 -424
rect 175 -526 209 -492
rect 271 -186 305 -152
rect 271 -254 305 -220
rect 271 -322 305 -288
rect 271 -390 305 -356
rect 271 -458 305 -424
rect 271 -526 305 -492
rect 367 -186 401 -152
rect 367 -254 401 -220
rect 367 -322 401 -288
rect 367 -390 401 -356
rect 367 -458 401 -424
rect 367 -526 401 -492
rect 463 -186 497 -152
rect 463 -254 497 -220
rect 463 -322 497 -288
rect 463 -390 497 -356
rect 463 -458 497 -424
rect 463 -526 497 -492
rect 559 -186 593 -152
rect 559 -254 593 -220
rect 559 -322 593 -288
rect 559 -390 593 -356
rect 559 -458 593 -424
rect 559 -526 593 -492
rect 655 -186 689 -152
rect 655 -254 689 -220
rect 655 -322 689 -288
rect 655 -390 689 -356
rect 655 -458 689 -424
rect 655 -526 689 -492
rect 751 -186 785 -152
rect 751 -254 785 -220
rect 751 -322 785 -288
rect 751 -390 785 -356
rect 751 -458 785 -424
rect 751 -526 785 -492
rect 847 -186 881 -152
rect 847 -254 881 -220
rect 847 -322 881 -288
rect 847 -390 881 -356
rect 847 -458 881 -424
rect 847 -526 881 -492
<< nsubdiff >>
rect -995 709 -867 743
rect -833 709 -799 743
rect -765 709 -731 743
rect -697 709 -663 743
rect -629 709 -595 743
rect -561 709 -527 743
rect -493 709 -459 743
rect -425 709 -391 743
rect -357 709 -323 743
rect -289 709 -255 743
rect -221 709 -187 743
rect -153 709 -119 743
rect -85 709 -51 743
rect -17 709 17 743
rect 51 709 85 743
rect 119 709 153 743
rect 187 709 221 743
rect 255 709 289 743
rect 323 709 357 743
rect 391 709 425 743
rect 459 709 493 743
rect 527 709 561 743
rect 595 709 629 743
rect 663 709 697 743
rect 731 709 765 743
rect 799 709 833 743
rect 867 709 995 743
rect -995 629 -961 709
rect -995 561 -961 595
rect 961 629 995 709
rect 961 561 995 595
rect -995 493 -961 527
rect -995 425 -961 459
rect -995 357 -961 391
rect -995 289 -961 323
rect -995 221 -961 255
rect -995 153 -961 187
rect -995 85 -961 119
rect 961 493 995 527
rect 961 425 995 459
rect 961 357 995 391
rect 961 289 995 323
rect 961 221 995 255
rect 961 153 995 187
rect -995 17 -961 51
rect 961 85 995 119
rect -995 -51 -961 -17
rect 961 17 995 51
rect -995 -119 -961 -85
rect 961 -51 995 -17
rect -995 -187 -961 -153
rect -995 -255 -961 -221
rect -995 -323 -961 -289
rect -995 -391 -961 -357
rect -995 -459 -961 -425
rect -995 -527 -961 -493
rect 961 -119 995 -85
rect 961 -187 995 -153
rect 961 -255 995 -221
rect 961 -323 995 -289
rect 961 -391 995 -357
rect 961 -459 995 -425
rect 961 -527 995 -493
rect -995 -595 -961 -561
rect -995 -709 -961 -629
rect 961 -595 995 -561
rect 961 -709 995 -629
rect -995 -743 -867 -709
rect -833 -743 -799 -709
rect -765 -743 -731 -709
rect -697 -743 -663 -709
rect -629 -743 -595 -709
rect -561 -743 -527 -709
rect -493 -743 -459 -709
rect -425 -743 -391 -709
rect -357 -743 -323 -709
rect -289 -743 -255 -709
rect -221 -743 -187 -709
rect -153 -743 -119 -709
rect -85 -743 -51 -709
rect -17 -743 17 -709
rect 51 -743 85 -709
rect 119 -743 153 -709
rect 187 -743 221 -709
rect 255 -743 289 -709
rect 323 -743 357 -709
rect 391 -743 425 -709
rect 459 -743 493 -709
rect 527 -743 561 -709
rect 595 -743 629 -709
rect 663 -743 697 -709
rect 731 -743 765 -709
rect 799 -743 833 -709
rect 867 -743 995 -709
<< nsubdiffcont >>
rect -867 709 -833 743
rect -799 709 -765 743
rect -731 709 -697 743
rect -663 709 -629 743
rect -595 709 -561 743
rect -527 709 -493 743
rect -459 709 -425 743
rect -391 709 -357 743
rect -323 709 -289 743
rect -255 709 -221 743
rect -187 709 -153 743
rect -119 709 -85 743
rect -51 709 -17 743
rect 17 709 51 743
rect 85 709 119 743
rect 153 709 187 743
rect 221 709 255 743
rect 289 709 323 743
rect 357 709 391 743
rect 425 709 459 743
rect 493 709 527 743
rect 561 709 595 743
rect 629 709 663 743
rect 697 709 731 743
rect 765 709 799 743
rect 833 709 867 743
rect -995 595 -961 629
rect 961 595 995 629
rect -995 527 -961 561
rect -995 459 -961 493
rect -995 391 -961 425
rect -995 323 -961 357
rect -995 255 -961 289
rect -995 187 -961 221
rect -995 119 -961 153
rect 961 527 995 561
rect 961 459 995 493
rect 961 391 995 425
rect 961 323 995 357
rect 961 255 995 289
rect 961 187 995 221
rect 961 119 995 153
rect -995 51 -961 85
rect 961 51 995 85
rect -995 -17 -961 17
rect 961 -17 995 17
rect -995 -85 -961 -51
rect 961 -85 995 -51
rect -995 -153 -961 -119
rect -995 -221 -961 -187
rect -995 -289 -961 -255
rect -995 -357 -961 -323
rect -995 -425 -961 -391
rect -995 -493 -961 -459
rect -995 -561 -961 -527
rect 961 -153 995 -119
rect 961 -221 995 -187
rect 961 -289 995 -255
rect 961 -357 995 -323
rect 961 -425 995 -391
rect 961 -493 995 -459
rect 961 -561 995 -527
rect -995 -629 -961 -595
rect 961 -629 995 -595
rect -867 -743 -833 -709
rect -799 -743 -765 -709
rect -731 -743 -697 -709
rect -663 -743 -629 -709
rect -595 -743 -561 -709
rect -527 -743 -493 -709
rect -459 -743 -425 -709
rect -391 -743 -357 -709
rect -323 -743 -289 -709
rect -255 -743 -221 -709
rect -187 -743 -153 -709
rect -119 -743 -85 -709
rect -51 -743 -17 -709
rect 17 -743 51 -709
rect 85 -743 119 -709
rect 153 -743 187 -709
rect 221 -743 255 -709
rect 289 -743 323 -709
rect 357 -743 391 -709
rect 425 -743 459 -709
rect 493 -743 527 -709
rect 561 -743 595 -709
rect 629 -743 663 -709
rect 697 -743 731 -709
rect 765 -743 799 -709
rect 833 -743 867 -709
<< poly >>
rect -849 641 -783 657
rect -849 607 -833 641
rect -799 607 -783 641
rect -849 591 -783 607
rect -657 641 -591 657
rect -657 607 -641 641
rect -607 607 -591 641
rect -657 591 -591 607
rect -465 641 -399 657
rect -465 607 -449 641
rect -415 607 -399 641
rect -465 591 -399 607
rect -273 641 -207 657
rect -273 607 -257 641
rect -223 607 -207 641
rect -273 591 -207 607
rect -81 641 -15 657
rect -81 607 -65 641
rect -31 607 -15 641
rect -81 591 -15 607
rect 111 641 177 657
rect 111 607 127 641
rect 161 607 177 641
rect 111 591 177 607
rect 303 641 369 657
rect 303 607 319 641
rect 353 607 369 641
rect 303 591 369 607
rect 495 641 561 657
rect 495 607 511 641
rect 545 607 561 641
rect 495 591 561 607
rect 687 641 753 657
rect 687 607 703 641
rect 737 607 753 641
rect 687 591 753 607
rect -831 560 -801 591
rect -735 560 -705 586
rect -639 560 -609 591
rect -543 560 -513 586
rect -447 560 -417 591
rect -351 560 -321 586
rect -255 560 -225 591
rect -159 560 -129 586
rect -63 560 -33 591
rect 33 560 63 586
rect 129 560 159 591
rect 225 560 255 586
rect 321 560 351 591
rect 417 560 447 586
rect 513 560 543 591
rect 609 560 639 586
rect 705 560 735 591
rect 801 560 831 586
rect -831 92 -801 118
rect -735 87 -705 118
rect -639 92 -609 118
rect -543 87 -513 118
rect -447 92 -417 118
rect -351 87 -321 118
rect -255 92 -225 118
rect -159 87 -129 118
rect -63 92 -33 118
rect 33 87 63 118
rect 129 92 159 118
rect 225 87 255 118
rect 321 92 351 118
rect 417 87 447 118
rect 513 92 543 118
rect 609 87 639 118
rect 705 92 735 118
rect 801 87 831 118
rect -753 71 -687 87
rect -753 37 -737 71
rect -703 37 -687 71
rect -753 21 -687 37
rect -561 71 -495 87
rect -561 37 -545 71
rect -511 37 -495 71
rect -561 21 -495 37
rect -369 71 -303 87
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect 591 71 657 87
rect 591 37 607 71
rect 641 37 657 71
rect 591 21 657 37
rect 783 71 849 87
rect 783 37 799 71
rect 833 37 849 71
rect 783 21 849 37
rect -753 -37 -687 -21
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -753 -87 -687 -71
rect -561 -37 -495 -21
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -561 -87 -495 -71
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 399 -87 465 -71
rect 591 -37 657 -21
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 591 -87 657 -71
rect 783 -37 849 -21
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 783 -87 849 -71
rect -831 -118 -801 -92
rect -735 -118 -705 -87
rect -639 -118 -609 -92
rect -543 -118 -513 -87
rect -447 -118 -417 -92
rect -351 -118 -321 -87
rect -255 -118 -225 -92
rect -159 -118 -129 -87
rect -63 -118 -33 -92
rect 33 -118 63 -87
rect 129 -118 159 -92
rect 225 -118 255 -87
rect 321 -118 351 -92
rect 417 -118 447 -87
rect 513 -118 543 -92
rect 609 -118 639 -87
rect 705 -118 735 -92
rect 801 -118 831 -87
rect -831 -591 -801 -560
rect -735 -586 -705 -560
rect -639 -591 -609 -560
rect -543 -586 -513 -560
rect -447 -591 -417 -560
rect -351 -586 -321 -560
rect -255 -591 -225 -560
rect -159 -586 -129 -560
rect -63 -591 -33 -560
rect 33 -586 63 -560
rect 129 -591 159 -560
rect 225 -586 255 -560
rect 321 -591 351 -560
rect 417 -586 447 -560
rect 513 -591 543 -560
rect 609 -586 639 -560
rect 705 -591 735 -560
rect 801 -586 831 -560
rect -849 -607 -783 -591
rect -849 -641 -833 -607
rect -799 -641 -783 -607
rect -849 -657 -783 -641
rect -657 -607 -591 -591
rect -657 -641 -641 -607
rect -607 -641 -591 -607
rect -657 -657 -591 -641
rect -465 -607 -399 -591
rect -465 -641 -449 -607
rect -415 -641 -399 -607
rect -465 -657 -399 -641
rect -273 -607 -207 -591
rect -273 -641 -257 -607
rect -223 -641 -207 -607
rect -273 -657 -207 -641
rect -81 -607 -15 -591
rect -81 -641 -65 -607
rect -31 -641 -15 -607
rect -81 -657 -15 -641
rect 111 -607 177 -591
rect 111 -641 127 -607
rect 161 -641 177 -607
rect 111 -657 177 -641
rect 303 -607 369 -591
rect 303 -641 319 -607
rect 353 -641 369 -607
rect 303 -657 369 -641
rect 495 -607 561 -591
rect 495 -641 511 -607
rect 545 -641 561 -607
rect 495 -657 561 -641
rect 687 -607 753 -591
rect 687 -641 703 -607
rect 737 -641 753 -607
rect 687 -657 753 -641
<< polycont >>
rect -833 607 -799 641
rect -641 607 -607 641
rect -449 607 -415 641
rect -257 607 -223 641
rect -65 607 -31 641
rect 127 607 161 641
rect 319 607 353 641
rect 511 607 545 641
rect 703 607 737 641
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect -833 -641 -799 -607
rect -641 -641 -607 -607
rect -449 -641 -415 -607
rect -257 -641 -223 -607
rect -65 -641 -31 -607
rect 127 -641 161 -607
rect 319 -641 353 -607
rect 511 -641 545 -607
rect 703 -641 737 -607
<< locali >>
rect -995 709 -867 743
rect -833 709 -799 743
rect -765 709 -731 743
rect -697 709 -663 743
rect -629 709 -595 743
rect -561 709 -527 743
rect -493 709 -459 743
rect -425 709 -391 743
rect -357 709 -323 743
rect -289 709 -255 743
rect -221 709 -187 743
rect -153 709 -119 743
rect -85 709 -51 743
rect -17 709 17 743
rect 51 709 85 743
rect 119 709 153 743
rect 187 709 221 743
rect 255 709 289 743
rect 323 709 357 743
rect 391 709 425 743
rect 459 709 493 743
rect 527 709 561 743
rect 595 709 629 743
rect 663 709 697 743
rect 731 709 765 743
rect 799 709 833 743
rect 867 709 995 743
rect -995 629 -961 709
rect -849 607 -833 641
rect -799 607 -783 641
rect -657 607 -641 641
rect -607 607 -591 641
rect -465 607 -449 641
rect -415 607 -399 641
rect -273 607 -257 641
rect -223 607 -207 641
rect -81 607 -65 641
rect -31 607 -15 641
rect 111 607 127 641
rect 161 607 177 641
rect 303 607 319 641
rect 353 607 369 641
rect 495 607 511 641
rect 545 607 561 641
rect 687 607 703 641
rect 737 607 753 641
rect 961 629 995 709
rect -995 561 -961 595
rect -995 493 -961 527
rect -995 425 -961 459
rect -995 357 -961 391
rect -995 289 -961 323
rect -995 221 -961 255
rect -995 153 -961 187
rect -995 85 -961 119
rect -881 536 -847 564
rect -881 464 -847 492
rect -881 392 -847 424
rect -881 322 -847 356
rect -881 254 -847 286
rect -881 186 -847 214
rect -881 114 -847 142
rect -785 536 -751 564
rect -785 464 -751 492
rect -785 392 -751 424
rect -785 322 -751 356
rect -785 254 -751 286
rect -785 186 -751 214
rect -785 114 -751 142
rect -689 536 -655 564
rect -689 464 -655 492
rect -689 392 -655 424
rect -689 322 -655 356
rect -689 254 -655 286
rect -689 186 -655 214
rect -689 114 -655 142
rect -593 536 -559 564
rect -593 464 -559 492
rect -593 392 -559 424
rect -593 322 -559 356
rect -593 254 -559 286
rect -593 186 -559 214
rect -593 114 -559 142
rect -497 536 -463 564
rect -497 464 -463 492
rect -497 392 -463 424
rect -497 322 -463 356
rect -497 254 -463 286
rect -497 186 -463 214
rect -497 114 -463 142
rect -401 536 -367 564
rect -401 464 -367 492
rect -401 392 -367 424
rect -401 322 -367 356
rect -401 254 -367 286
rect -401 186 -367 214
rect -401 114 -367 142
rect -305 536 -271 564
rect -305 464 -271 492
rect -305 392 -271 424
rect -305 322 -271 356
rect -305 254 -271 286
rect -305 186 -271 214
rect -305 114 -271 142
rect -209 536 -175 564
rect -209 464 -175 492
rect -209 392 -175 424
rect -209 322 -175 356
rect -209 254 -175 286
rect -209 186 -175 214
rect -209 114 -175 142
rect -113 536 -79 564
rect -113 464 -79 492
rect -113 392 -79 424
rect -113 322 -79 356
rect -113 254 -79 286
rect -113 186 -79 214
rect -113 114 -79 142
rect -17 536 17 564
rect -17 464 17 492
rect -17 392 17 424
rect -17 322 17 356
rect -17 254 17 286
rect -17 186 17 214
rect -17 114 17 142
rect 79 536 113 564
rect 79 464 113 492
rect 79 392 113 424
rect 79 322 113 356
rect 79 254 113 286
rect 79 186 113 214
rect 79 114 113 142
rect 175 536 209 564
rect 175 464 209 492
rect 175 392 209 424
rect 175 322 209 356
rect 175 254 209 286
rect 175 186 209 214
rect 175 114 209 142
rect 271 536 305 564
rect 271 464 305 492
rect 271 392 305 424
rect 271 322 305 356
rect 271 254 305 286
rect 271 186 305 214
rect 271 114 305 142
rect 367 536 401 564
rect 367 464 401 492
rect 367 392 401 424
rect 367 322 401 356
rect 367 254 401 286
rect 367 186 401 214
rect 367 114 401 142
rect 463 536 497 564
rect 463 464 497 492
rect 463 392 497 424
rect 463 322 497 356
rect 463 254 497 286
rect 463 186 497 214
rect 463 114 497 142
rect 559 536 593 564
rect 559 464 593 492
rect 559 392 593 424
rect 559 322 593 356
rect 559 254 593 286
rect 559 186 593 214
rect 559 114 593 142
rect 655 536 689 564
rect 655 464 689 492
rect 655 392 689 424
rect 655 322 689 356
rect 655 254 689 286
rect 655 186 689 214
rect 655 114 689 142
rect 751 536 785 564
rect 751 464 785 492
rect 751 392 785 424
rect 751 322 785 356
rect 751 254 785 286
rect 751 186 785 214
rect 751 114 785 142
rect 847 536 881 564
rect 847 464 881 492
rect 847 392 881 424
rect 847 322 881 356
rect 847 254 881 286
rect 847 186 881 214
rect 847 114 881 142
rect 961 561 995 595
rect 961 493 995 527
rect 961 425 995 459
rect 961 357 995 391
rect 961 289 995 323
rect 961 221 995 255
rect 961 153 995 187
rect 961 85 995 119
rect -995 17 -961 51
rect -753 37 -737 71
rect -703 37 -687 71
rect -561 37 -545 71
rect -511 37 -495 71
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect 591 37 607 71
rect 641 37 657 71
rect 783 37 799 71
rect 833 37 849 71
rect -995 -51 -961 -17
rect 961 17 995 51
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 961 -51 995 -17
rect -995 -119 -961 -85
rect -995 -187 -961 -153
rect -995 -255 -961 -221
rect -995 -323 -961 -289
rect -995 -391 -961 -357
rect -995 -459 -961 -425
rect -995 -527 -961 -493
rect -995 -595 -961 -561
rect -881 -142 -847 -114
rect -881 -214 -847 -186
rect -881 -286 -847 -254
rect -881 -356 -847 -322
rect -881 -424 -847 -392
rect -881 -492 -847 -464
rect -881 -564 -847 -536
rect -785 -142 -751 -114
rect -785 -214 -751 -186
rect -785 -286 -751 -254
rect -785 -356 -751 -322
rect -785 -424 -751 -392
rect -785 -492 -751 -464
rect -785 -564 -751 -536
rect -689 -142 -655 -114
rect -689 -214 -655 -186
rect -689 -286 -655 -254
rect -689 -356 -655 -322
rect -689 -424 -655 -392
rect -689 -492 -655 -464
rect -689 -564 -655 -536
rect -593 -142 -559 -114
rect -593 -214 -559 -186
rect -593 -286 -559 -254
rect -593 -356 -559 -322
rect -593 -424 -559 -392
rect -593 -492 -559 -464
rect -593 -564 -559 -536
rect -497 -142 -463 -114
rect -497 -214 -463 -186
rect -497 -286 -463 -254
rect -497 -356 -463 -322
rect -497 -424 -463 -392
rect -497 -492 -463 -464
rect -497 -564 -463 -536
rect -401 -142 -367 -114
rect -401 -214 -367 -186
rect -401 -286 -367 -254
rect -401 -356 -367 -322
rect -401 -424 -367 -392
rect -401 -492 -367 -464
rect -401 -564 -367 -536
rect -305 -142 -271 -114
rect -305 -214 -271 -186
rect -305 -286 -271 -254
rect -305 -356 -271 -322
rect -305 -424 -271 -392
rect -305 -492 -271 -464
rect -305 -564 -271 -536
rect -209 -142 -175 -114
rect -209 -214 -175 -186
rect -209 -286 -175 -254
rect -209 -356 -175 -322
rect -209 -424 -175 -392
rect -209 -492 -175 -464
rect -209 -564 -175 -536
rect -113 -142 -79 -114
rect -113 -214 -79 -186
rect -113 -286 -79 -254
rect -113 -356 -79 -322
rect -113 -424 -79 -392
rect -113 -492 -79 -464
rect -113 -564 -79 -536
rect -17 -142 17 -114
rect -17 -214 17 -186
rect -17 -286 17 -254
rect -17 -356 17 -322
rect -17 -424 17 -392
rect -17 -492 17 -464
rect -17 -564 17 -536
rect 79 -142 113 -114
rect 79 -214 113 -186
rect 79 -286 113 -254
rect 79 -356 113 -322
rect 79 -424 113 -392
rect 79 -492 113 -464
rect 79 -564 113 -536
rect 175 -142 209 -114
rect 175 -214 209 -186
rect 175 -286 209 -254
rect 175 -356 209 -322
rect 175 -424 209 -392
rect 175 -492 209 -464
rect 175 -564 209 -536
rect 271 -142 305 -114
rect 271 -214 305 -186
rect 271 -286 305 -254
rect 271 -356 305 -322
rect 271 -424 305 -392
rect 271 -492 305 -464
rect 271 -564 305 -536
rect 367 -142 401 -114
rect 367 -214 401 -186
rect 367 -286 401 -254
rect 367 -356 401 -322
rect 367 -424 401 -392
rect 367 -492 401 -464
rect 367 -564 401 -536
rect 463 -142 497 -114
rect 463 -214 497 -186
rect 463 -286 497 -254
rect 463 -356 497 -322
rect 463 -424 497 -392
rect 463 -492 497 -464
rect 463 -564 497 -536
rect 559 -142 593 -114
rect 559 -214 593 -186
rect 559 -286 593 -254
rect 559 -356 593 -322
rect 559 -424 593 -392
rect 559 -492 593 -464
rect 559 -564 593 -536
rect 655 -142 689 -114
rect 655 -214 689 -186
rect 655 -286 689 -254
rect 655 -356 689 -322
rect 655 -424 689 -392
rect 655 -492 689 -464
rect 655 -564 689 -536
rect 751 -142 785 -114
rect 751 -214 785 -186
rect 751 -286 785 -254
rect 751 -356 785 -322
rect 751 -424 785 -392
rect 751 -492 785 -464
rect 751 -564 785 -536
rect 847 -142 881 -114
rect 847 -214 881 -186
rect 847 -286 881 -254
rect 847 -356 881 -322
rect 847 -424 881 -392
rect 847 -492 881 -464
rect 847 -564 881 -536
rect 961 -119 995 -85
rect 961 -187 995 -153
rect 961 -255 995 -221
rect 961 -323 995 -289
rect 961 -391 995 -357
rect 961 -459 995 -425
rect 961 -527 995 -493
rect 961 -595 995 -561
rect -995 -709 -961 -629
rect -849 -641 -833 -607
rect -799 -641 -783 -607
rect -657 -641 -641 -607
rect -607 -641 -591 -607
rect -465 -641 -449 -607
rect -415 -641 -399 -607
rect -273 -641 -257 -607
rect -223 -641 -207 -607
rect -81 -641 -65 -607
rect -31 -641 -15 -607
rect 111 -641 127 -607
rect 161 -641 177 -607
rect 303 -641 319 -607
rect 353 -641 369 -607
rect 495 -641 511 -607
rect 545 -641 561 -607
rect 687 -641 703 -607
rect 737 -641 753 -607
rect 961 -709 995 -629
rect -995 -743 -867 -709
rect -833 -743 -799 -709
rect -765 -743 -731 -709
rect -697 -743 -663 -709
rect -629 -743 -595 -709
rect -561 -743 -527 -709
rect -493 -743 -459 -709
rect -425 -743 -391 -709
rect -357 -743 -323 -709
rect -289 -743 -255 -709
rect -221 -743 -187 -709
rect -153 -743 -119 -709
rect -85 -743 -51 -709
rect -17 -743 17 -709
rect 51 -743 85 -709
rect 119 -743 153 -709
rect 187 -743 221 -709
rect 255 -743 289 -709
rect 323 -743 357 -709
rect 391 -743 425 -709
rect 459 -743 493 -709
rect 527 -743 561 -709
rect 595 -743 629 -709
rect 663 -743 697 -709
rect 731 -743 765 -709
rect 799 -743 833 -709
rect 867 -743 995 -709
<< viali >>
rect -833 607 -799 641
rect -641 607 -607 641
rect -449 607 -415 641
rect -257 607 -223 641
rect -65 607 -31 641
rect 127 607 161 641
rect 319 607 353 641
rect 511 607 545 641
rect 703 607 737 641
rect -881 526 -847 536
rect -881 502 -847 526
rect -881 458 -847 464
rect -881 430 -847 458
rect -881 390 -847 392
rect -881 358 -847 390
rect -881 288 -847 320
rect -881 286 -847 288
rect -881 220 -847 248
rect -881 214 -847 220
rect -881 152 -847 176
rect -881 142 -847 152
rect -785 526 -751 536
rect -785 502 -751 526
rect -785 458 -751 464
rect -785 430 -751 458
rect -785 390 -751 392
rect -785 358 -751 390
rect -785 288 -751 320
rect -785 286 -751 288
rect -785 220 -751 248
rect -785 214 -751 220
rect -785 152 -751 176
rect -785 142 -751 152
rect -689 526 -655 536
rect -689 502 -655 526
rect -689 458 -655 464
rect -689 430 -655 458
rect -689 390 -655 392
rect -689 358 -655 390
rect -689 288 -655 320
rect -689 286 -655 288
rect -689 220 -655 248
rect -689 214 -655 220
rect -689 152 -655 176
rect -689 142 -655 152
rect -593 526 -559 536
rect -593 502 -559 526
rect -593 458 -559 464
rect -593 430 -559 458
rect -593 390 -559 392
rect -593 358 -559 390
rect -593 288 -559 320
rect -593 286 -559 288
rect -593 220 -559 248
rect -593 214 -559 220
rect -593 152 -559 176
rect -593 142 -559 152
rect -497 526 -463 536
rect -497 502 -463 526
rect -497 458 -463 464
rect -497 430 -463 458
rect -497 390 -463 392
rect -497 358 -463 390
rect -497 288 -463 320
rect -497 286 -463 288
rect -497 220 -463 248
rect -497 214 -463 220
rect -497 152 -463 176
rect -497 142 -463 152
rect -401 526 -367 536
rect -401 502 -367 526
rect -401 458 -367 464
rect -401 430 -367 458
rect -401 390 -367 392
rect -401 358 -367 390
rect -401 288 -367 320
rect -401 286 -367 288
rect -401 220 -367 248
rect -401 214 -367 220
rect -401 152 -367 176
rect -401 142 -367 152
rect -305 526 -271 536
rect -305 502 -271 526
rect -305 458 -271 464
rect -305 430 -271 458
rect -305 390 -271 392
rect -305 358 -271 390
rect -305 288 -271 320
rect -305 286 -271 288
rect -305 220 -271 248
rect -305 214 -271 220
rect -305 152 -271 176
rect -305 142 -271 152
rect -209 526 -175 536
rect -209 502 -175 526
rect -209 458 -175 464
rect -209 430 -175 458
rect -209 390 -175 392
rect -209 358 -175 390
rect -209 288 -175 320
rect -209 286 -175 288
rect -209 220 -175 248
rect -209 214 -175 220
rect -209 152 -175 176
rect -209 142 -175 152
rect -113 526 -79 536
rect -113 502 -79 526
rect -113 458 -79 464
rect -113 430 -79 458
rect -113 390 -79 392
rect -113 358 -79 390
rect -113 288 -79 320
rect -113 286 -79 288
rect -113 220 -79 248
rect -113 214 -79 220
rect -113 152 -79 176
rect -113 142 -79 152
rect -17 526 17 536
rect -17 502 17 526
rect -17 458 17 464
rect -17 430 17 458
rect -17 390 17 392
rect -17 358 17 390
rect -17 288 17 320
rect -17 286 17 288
rect -17 220 17 248
rect -17 214 17 220
rect -17 152 17 176
rect -17 142 17 152
rect 79 526 113 536
rect 79 502 113 526
rect 79 458 113 464
rect 79 430 113 458
rect 79 390 113 392
rect 79 358 113 390
rect 79 288 113 320
rect 79 286 113 288
rect 79 220 113 248
rect 79 214 113 220
rect 79 152 113 176
rect 79 142 113 152
rect 175 526 209 536
rect 175 502 209 526
rect 175 458 209 464
rect 175 430 209 458
rect 175 390 209 392
rect 175 358 209 390
rect 175 288 209 320
rect 175 286 209 288
rect 175 220 209 248
rect 175 214 209 220
rect 175 152 209 176
rect 175 142 209 152
rect 271 526 305 536
rect 271 502 305 526
rect 271 458 305 464
rect 271 430 305 458
rect 271 390 305 392
rect 271 358 305 390
rect 271 288 305 320
rect 271 286 305 288
rect 271 220 305 248
rect 271 214 305 220
rect 271 152 305 176
rect 271 142 305 152
rect 367 526 401 536
rect 367 502 401 526
rect 367 458 401 464
rect 367 430 401 458
rect 367 390 401 392
rect 367 358 401 390
rect 367 288 401 320
rect 367 286 401 288
rect 367 220 401 248
rect 367 214 401 220
rect 367 152 401 176
rect 367 142 401 152
rect 463 526 497 536
rect 463 502 497 526
rect 463 458 497 464
rect 463 430 497 458
rect 463 390 497 392
rect 463 358 497 390
rect 463 288 497 320
rect 463 286 497 288
rect 463 220 497 248
rect 463 214 497 220
rect 463 152 497 176
rect 463 142 497 152
rect 559 526 593 536
rect 559 502 593 526
rect 559 458 593 464
rect 559 430 593 458
rect 559 390 593 392
rect 559 358 593 390
rect 559 288 593 320
rect 559 286 593 288
rect 559 220 593 248
rect 559 214 593 220
rect 559 152 593 176
rect 559 142 593 152
rect 655 526 689 536
rect 655 502 689 526
rect 655 458 689 464
rect 655 430 689 458
rect 655 390 689 392
rect 655 358 689 390
rect 655 288 689 320
rect 655 286 689 288
rect 655 220 689 248
rect 655 214 689 220
rect 655 152 689 176
rect 655 142 689 152
rect 751 526 785 536
rect 751 502 785 526
rect 751 458 785 464
rect 751 430 785 458
rect 751 390 785 392
rect 751 358 785 390
rect 751 288 785 320
rect 751 286 785 288
rect 751 220 785 248
rect 751 214 785 220
rect 751 152 785 176
rect 751 142 785 152
rect 847 526 881 536
rect 847 502 881 526
rect 847 458 881 464
rect 847 430 881 458
rect 847 390 881 392
rect 847 358 881 390
rect 847 288 881 320
rect 847 286 881 288
rect 847 220 881 248
rect 847 214 881 220
rect 847 152 881 176
rect 847 142 881 152
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect -881 -152 -847 -142
rect -881 -176 -847 -152
rect -881 -220 -847 -214
rect -881 -248 -847 -220
rect -881 -288 -847 -286
rect -881 -320 -847 -288
rect -881 -390 -847 -358
rect -881 -392 -847 -390
rect -881 -458 -847 -430
rect -881 -464 -847 -458
rect -881 -526 -847 -502
rect -881 -536 -847 -526
rect -785 -152 -751 -142
rect -785 -176 -751 -152
rect -785 -220 -751 -214
rect -785 -248 -751 -220
rect -785 -288 -751 -286
rect -785 -320 -751 -288
rect -785 -390 -751 -358
rect -785 -392 -751 -390
rect -785 -458 -751 -430
rect -785 -464 -751 -458
rect -785 -526 -751 -502
rect -785 -536 -751 -526
rect -689 -152 -655 -142
rect -689 -176 -655 -152
rect -689 -220 -655 -214
rect -689 -248 -655 -220
rect -689 -288 -655 -286
rect -689 -320 -655 -288
rect -689 -390 -655 -358
rect -689 -392 -655 -390
rect -689 -458 -655 -430
rect -689 -464 -655 -458
rect -689 -526 -655 -502
rect -689 -536 -655 -526
rect -593 -152 -559 -142
rect -593 -176 -559 -152
rect -593 -220 -559 -214
rect -593 -248 -559 -220
rect -593 -288 -559 -286
rect -593 -320 -559 -288
rect -593 -390 -559 -358
rect -593 -392 -559 -390
rect -593 -458 -559 -430
rect -593 -464 -559 -458
rect -593 -526 -559 -502
rect -593 -536 -559 -526
rect -497 -152 -463 -142
rect -497 -176 -463 -152
rect -497 -220 -463 -214
rect -497 -248 -463 -220
rect -497 -288 -463 -286
rect -497 -320 -463 -288
rect -497 -390 -463 -358
rect -497 -392 -463 -390
rect -497 -458 -463 -430
rect -497 -464 -463 -458
rect -497 -526 -463 -502
rect -497 -536 -463 -526
rect -401 -152 -367 -142
rect -401 -176 -367 -152
rect -401 -220 -367 -214
rect -401 -248 -367 -220
rect -401 -288 -367 -286
rect -401 -320 -367 -288
rect -401 -390 -367 -358
rect -401 -392 -367 -390
rect -401 -458 -367 -430
rect -401 -464 -367 -458
rect -401 -526 -367 -502
rect -401 -536 -367 -526
rect -305 -152 -271 -142
rect -305 -176 -271 -152
rect -305 -220 -271 -214
rect -305 -248 -271 -220
rect -305 -288 -271 -286
rect -305 -320 -271 -288
rect -305 -390 -271 -358
rect -305 -392 -271 -390
rect -305 -458 -271 -430
rect -305 -464 -271 -458
rect -305 -526 -271 -502
rect -305 -536 -271 -526
rect -209 -152 -175 -142
rect -209 -176 -175 -152
rect -209 -220 -175 -214
rect -209 -248 -175 -220
rect -209 -288 -175 -286
rect -209 -320 -175 -288
rect -209 -390 -175 -358
rect -209 -392 -175 -390
rect -209 -458 -175 -430
rect -209 -464 -175 -458
rect -209 -526 -175 -502
rect -209 -536 -175 -526
rect -113 -152 -79 -142
rect -113 -176 -79 -152
rect -113 -220 -79 -214
rect -113 -248 -79 -220
rect -113 -288 -79 -286
rect -113 -320 -79 -288
rect -113 -390 -79 -358
rect -113 -392 -79 -390
rect -113 -458 -79 -430
rect -113 -464 -79 -458
rect -113 -526 -79 -502
rect -113 -536 -79 -526
rect -17 -152 17 -142
rect -17 -176 17 -152
rect -17 -220 17 -214
rect -17 -248 17 -220
rect -17 -288 17 -286
rect -17 -320 17 -288
rect -17 -390 17 -358
rect -17 -392 17 -390
rect -17 -458 17 -430
rect -17 -464 17 -458
rect -17 -526 17 -502
rect -17 -536 17 -526
rect 79 -152 113 -142
rect 79 -176 113 -152
rect 79 -220 113 -214
rect 79 -248 113 -220
rect 79 -288 113 -286
rect 79 -320 113 -288
rect 79 -390 113 -358
rect 79 -392 113 -390
rect 79 -458 113 -430
rect 79 -464 113 -458
rect 79 -526 113 -502
rect 79 -536 113 -526
rect 175 -152 209 -142
rect 175 -176 209 -152
rect 175 -220 209 -214
rect 175 -248 209 -220
rect 175 -288 209 -286
rect 175 -320 209 -288
rect 175 -390 209 -358
rect 175 -392 209 -390
rect 175 -458 209 -430
rect 175 -464 209 -458
rect 175 -526 209 -502
rect 175 -536 209 -526
rect 271 -152 305 -142
rect 271 -176 305 -152
rect 271 -220 305 -214
rect 271 -248 305 -220
rect 271 -288 305 -286
rect 271 -320 305 -288
rect 271 -390 305 -358
rect 271 -392 305 -390
rect 271 -458 305 -430
rect 271 -464 305 -458
rect 271 -526 305 -502
rect 271 -536 305 -526
rect 367 -152 401 -142
rect 367 -176 401 -152
rect 367 -220 401 -214
rect 367 -248 401 -220
rect 367 -288 401 -286
rect 367 -320 401 -288
rect 367 -390 401 -358
rect 367 -392 401 -390
rect 367 -458 401 -430
rect 367 -464 401 -458
rect 367 -526 401 -502
rect 367 -536 401 -526
rect 463 -152 497 -142
rect 463 -176 497 -152
rect 463 -220 497 -214
rect 463 -248 497 -220
rect 463 -288 497 -286
rect 463 -320 497 -288
rect 463 -390 497 -358
rect 463 -392 497 -390
rect 463 -458 497 -430
rect 463 -464 497 -458
rect 463 -526 497 -502
rect 463 -536 497 -526
rect 559 -152 593 -142
rect 559 -176 593 -152
rect 559 -220 593 -214
rect 559 -248 593 -220
rect 559 -288 593 -286
rect 559 -320 593 -288
rect 559 -390 593 -358
rect 559 -392 593 -390
rect 559 -458 593 -430
rect 559 -464 593 -458
rect 559 -526 593 -502
rect 559 -536 593 -526
rect 655 -152 689 -142
rect 655 -176 689 -152
rect 655 -220 689 -214
rect 655 -248 689 -220
rect 655 -288 689 -286
rect 655 -320 689 -288
rect 655 -390 689 -358
rect 655 -392 689 -390
rect 655 -458 689 -430
rect 655 -464 689 -458
rect 655 -526 689 -502
rect 655 -536 689 -526
rect 751 -152 785 -142
rect 751 -176 785 -152
rect 751 -220 785 -214
rect 751 -248 785 -220
rect 751 -288 785 -286
rect 751 -320 785 -288
rect 751 -390 785 -358
rect 751 -392 785 -390
rect 751 -458 785 -430
rect 751 -464 785 -458
rect 751 -526 785 -502
rect 751 -536 785 -526
rect 847 -152 881 -142
rect 847 -176 881 -152
rect 847 -220 881 -214
rect 847 -248 881 -220
rect 847 -288 881 -286
rect 847 -320 881 -288
rect 847 -390 881 -358
rect 847 -392 881 -390
rect 847 -458 881 -430
rect 847 -464 881 -458
rect 847 -526 881 -502
rect 847 -536 881 -526
rect -833 -641 -799 -607
rect -641 -641 -607 -607
rect -449 -641 -415 -607
rect -257 -641 -223 -607
rect -65 -641 -31 -607
rect 127 -641 161 -607
rect 319 -641 353 -607
rect 511 -641 545 -607
rect 703 -641 737 -607
<< metal1 >>
rect -845 641 -787 647
rect -845 607 -833 641
rect -799 607 -787 641
rect -845 601 -787 607
rect -653 641 -595 647
rect -653 607 -641 641
rect -607 607 -595 641
rect -653 601 -595 607
rect -461 641 -403 647
rect -461 607 -449 641
rect -415 607 -403 641
rect -461 601 -403 607
rect -269 641 -211 647
rect -269 607 -257 641
rect -223 607 -211 641
rect -269 601 -211 607
rect -77 641 -19 647
rect -77 607 -65 641
rect -31 607 -19 641
rect -77 601 -19 607
rect 115 641 173 647
rect 115 607 127 641
rect 161 607 173 641
rect 115 601 173 607
rect 307 641 365 647
rect 307 607 319 641
rect 353 607 365 641
rect 307 601 365 607
rect 499 641 557 647
rect 499 607 511 641
rect 545 607 557 641
rect 499 601 557 607
rect 691 641 749 647
rect 691 607 703 641
rect 737 607 749 641
rect 691 601 749 607
rect -887 536 -841 560
rect -887 502 -881 536
rect -847 502 -841 536
rect -887 464 -841 502
rect -887 430 -881 464
rect -847 430 -841 464
rect -887 392 -841 430
rect -887 358 -881 392
rect -847 358 -841 392
rect -887 320 -841 358
rect -887 286 -881 320
rect -847 286 -841 320
rect -887 248 -841 286
rect -887 214 -881 248
rect -847 214 -841 248
rect -887 176 -841 214
rect -887 142 -881 176
rect -847 142 -841 176
rect -887 118 -841 142
rect -791 536 -745 560
rect -791 502 -785 536
rect -751 502 -745 536
rect -791 464 -745 502
rect -791 430 -785 464
rect -751 430 -745 464
rect -791 392 -745 430
rect -791 358 -785 392
rect -751 358 -745 392
rect -791 320 -745 358
rect -791 286 -785 320
rect -751 286 -745 320
rect -791 248 -745 286
rect -791 214 -785 248
rect -751 214 -745 248
rect -791 176 -745 214
rect -791 142 -785 176
rect -751 142 -745 176
rect -791 118 -745 142
rect -695 536 -649 560
rect -695 502 -689 536
rect -655 502 -649 536
rect -695 464 -649 502
rect -695 430 -689 464
rect -655 430 -649 464
rect -695 392 -649 430
rect -695 358 -689 392
rect -655 358 -649 392
rect -695 320 -649 358
rect -695 286 -689 320
rect -655 286 -649 320
rect -695 248 -649 286
rect -695 214 -689 248
rect -655 214 -649 248
rect -695 176 -649 214
rect -695 142 -689 176
rect -655 142 -649 176
rect -695 118 -649 142
rect -599 536 -553 560
rect -599 502 -593 536
rect -559 502 -553 536
rect -599 464 -553 502
rect -599 430 -593 464
rect -559 430 -553 464
rect -599 392 -553 430
rect -599 358 -593 392
rect -559 358 -553 392
rect -599 320 -553 358
rect -599 286 -593 320
rect -559 286 -553 320
rect -599 248 -553 286
rect -599 214 -593 248
rect -559 214 -553 248
rect -599 176 -553 214
rect -599 142 -593 176
rect -559 142 -553 176
rect -599 118 -553 142
rect -503 536 -457 560
rect -503 502 -497 536
rect -463 502 -457 536
rect -503 464 -457 502
rect -503 430 -497 464
rect -463 430 -457 464
rect -503 392 -457 430
rect -503 358 -497 392
rect -463 358 -457 392
rect -503 320 -457 358
rect -503 286 -497 320
rect -463 286 -457 320
rect -503 248 -457 286
rect -503 214 -497 248
rect -463 214 -457 248
rect -503 176 -457 214
rect -503 142 -497 176
rect -463 142 -457 176
rect -503 118 -457 142
rect -407 536 -361 560
rect -407 502 -401 536
rect -367 502 -361 536
rect -407 464 -361 502
rect -407 430 -401 464
rect -367 430 -361 464
rect -407 392 -361 430
rect -407 358 -401 392
rect -367 358 -361 392
rect -407 320 -361 358
rect -407 286 -401 320
rect -367 286 -361 320
rect -407 248 -361 286
rect -407 214 -401 248
rect -367 214 -361 248
rect -407 176 -361 214
rect -407 142 -401 176
rect -367 142 -361 176
rect -407 118 -361 142
rect -311 536 -265 560
rect -311 502 -305 536
rect -271 502 -265 536
rect -311 464 -265 502
rect -311 430 -305 464
rect -271 430 -265 464
rect -311 392 -265 430
rect -311 358 -305 392
rect -271 358 -265 392
rect -311 320 -265 358
rect -311 286 -305 320
rect -271 286 -265 320
rect -311 248 -265 286
rect -311 214 -305 248
rect -271 214 -265 248
rect -311 176 -265 214
rect -311 142 -305 176
rect -271 142 -265 176
rect -311 118 -265 142
rect -215 536 -169 560
rect -215 502 -209 536
rect -175 502 -169 536
rect -215 464 -169 502
rect -215 430 -209 464
rect -175 430 -169 464
rect -215 392 -169 430
rect -215 358 -209 392
rect -175 358 -169 392
rect -215 320 -169 358
rect -215 286 -209 320
rect -175 286 -169 320
rect -215 248 -169 286
rect -215 214 -209 248
rect -175 214 -169 248
rect -215 176 -169 214
rect -215 142 -209 176
rect -175 142 -169 176
rect -215 118 -169 142
rect -119 536 -73 560
rect -119 502 -113 536
rect -79 502 -73 536
rect -119 464 -73 502
rect -119 430 -113 464
rect -79 430 -73 464
rect -119 392 -73 430
rect -119 358 -113 392
rect -79 358 -73 392
rect -119 320 -73 358
rect -119 286 -113 320
rect -79 286 -73 320
rect -119 248 -73 286
rect -119 214 -113 248
rect -79 214 -73 248
rect -119 176 -73 214
rect -119 142 -113 176
rect -79 142 -73 176
rect -119 118 -73 142
rect -23 536 23 560
rect -23 502 -17 536
rect 17 502 23 536
rect -23 464 23 502
rect -23 430 -17 464
rect 17 430 23 464
rect -23 392 23 430
rect -23 358 -17 392
rect 17 358 23 392
rect -23 320 23 358
rect -23 286 -17 320
rect 17 286 23 320
rect -23 248 23 286
rect -23 214 -17 248
rect 17 214 23 248
rect -23 176 23 214
rect -23 142 -17 176
rect 17 142 23 176
rect -23 118 23 142
rect 73 536 119 560
rect 73 502 79 536
rect 113 502 119 536
rect 73 464 119 502
rect 73 430 79 464
rect 113 430 119 464
rect 73 392 119 430
rect 73 358 79 392
rect 113 358 119 392
rect 73 320 119 358
rect 73 286 79 320
rect 113 286 119 320
rect 73 248 119 286
rect 73 214 79 248
rect 113 214 119 248
rect 73 176 119 214
rect 73 142 79 176
rect 113 142 119 176
rect 73 118 119 142
rect 169 536 215 560
rect 169 502 175 536
rect 209 502 215 536
rect 169 464 215 502
rect 169 430 175 464
rect 209 430 215 464
rect 169 392 215 430
rect 169 358 175 392
rect 209 358 215 392
rect 169 320 215 358
rect 169 286 175 320
rect 209 286 215 320
rect 169 248 215 286
rect 169 214 175 248
rect 209 214 215 248
rect 169 176 215 214
rect 169 142 175 176
rect 209 142 215 176
rect 169 118 215 142
rect 265 536 311 560
rect 265 502 271 536
rect 305 502 311 536
rect 265 464 311 502
rect 265 430 271 464
rect 305 430 311 464
rect 265 392 311 430
rect 265 358 271 392
rect 305 358 311 392
rect 265 320 311 358
rect 265 286 271 320
rect 305 286 311 320
rect 265 248 311 286
rect 265 214 271 248
rect 305 214 311 248
rect 265 176 311 214
rect 265 142 271 176
rect 305 142 311 176
rect 265 118 311 142
rect 361 536 407 560
rect 361 502 367 536
rect 401 502 407 536
rect 361 464 407 502
rect 361 430 367 464
rect 401 430 407 464
rect 361 392 407 430
rect 361 358 367 392
rect 401 358 407 392
rect 361 320 407 358
rect 361 286 367 320
rect 401 286 407 320
rect 361 248 407 286
rect 361 214 367 248
rect 401 214 407 248
rect 361 176 407 214
rect 361 142 367 176
rect 401 142 407 176
rect 361 118 407 142
rect 457 536 503 560
rect 457 502 463 536
rect 497 502 503 536
rect 457 464 503 502
rect 457 430 463 464
rect 497 430 503 464
rect 457 392 503 430
rect 457 358 463 392
rect 497 358 503 392
rect 457 320 503 358
rect 457 286 463 320
rect 497 286 503 320
rect 457 248 503 286
rect 457 214 463 248
rect 497 214 503 248
rect 457 176 503 214
rect 457 142 463 176
rect 497 142 503 176
rect 457 118 503 142
rect 553 536 599 560
rect 553 502 559 536
rect 593 502 599 536
rect 553 464 599 502
rect 553 430 559 464
rect 593 430 599 464
rect 553 392 599 430
rect 553 358 559 392
rect 593 358 599 392
rect 553 320 599 358
rect 553 286 559 320
rect 593 286 599 320
rect 553 248 599 286
rect 553 214 559 248
rect 593 214 599 248
rect 553 176 599 214
rect 553 142 559 176
rect 593 142 599 176
rect 553 118 599 142
rect 649 536 695 560
rect 649 502 655 536
rect 689 502 695 536
rect 649 464 695 502
rect 649 430 655 464
rect 689 430 695 464
rect 649 392 695 430
rect 649 358 655 392
rect 689 358 695 392
rect 649 320 695 358
rect 649 286 655 320
rect 689 286 695 320
rect 649 248 695 286
rect 649 214 655 248
rect 689 214 695 248
rect 649 176 695 214
rect 649 142 655 176
rect 689 142 695 176
rect 649 118 695 142
rect 745 536 791 560
rect 745 502 751 536
rect 785 502 791 536
rect 745 464 791 502
rect 745 430 751 464
rect 785 430 791 464
rect 745 392 791 430
rect 745 358 751 392
rect 785 358 791 392
rect 745 320 791 358
rect 745 286 751 320
rect 785 286 791 320
rect 745 248 791 286
rect 745 214 751 248
rect 785 214 791 248
rect 745 176 791 214
rect 745 142 751 176
rect 785 142 791 176
rect 745 118 791 142
rect 841 536 887 560
rect 841 502 847 536
rect 881 502 887 536
rect 841 464 887 502
rect 841 430 847 464
rect 881 430 887 464
rect 841 392 887 430
rect 841 358 847 392
rect 881 358 887 392
rect 841 320 887 358
rect 841 286 847 320
rect 881 286 887 320
rect 841 248 887 286
rect 841 214 847 248
rect 881 214 887 248
rect 841 176 887 214
rect 841 142 847 176
rect 881 142 887 176
rect 841 118 887 142
rect -749 71 -691 77
rect -749 37 -737 71
rect -703 37 -691 71
rect -749 31 -691 37
rect -557 71 -499 77
rect -557 37 -545 71
rect -511 37 -499 71
rect -557 31 -499 37
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect 595 71 653 77
rect 595 37 607 71
rect 641 37 653 71
rect 595 31 653 37
rect 787 71 845 77
rect 787 37 799 71
rect 833 37 845 71
rect 787 31 845 37
rect -749 -37 -691 -31
rect -749 -71 -737 -37
rect -703 -71 -691 -37
rect -749 -77 -691 -71
rect -557 -37 -499 -31
rect -557 -71 -545 -37
rect -511 -71 -499 -37
rect -557 -77 -499 -71
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect 595 -37 653 -31
rect 595 -71 607 -37
rect 641 -71 653 -37
rect 595 -77 653 -71
rect 787 -37 845 -31
rect 787 -71 799 -37
rect 833 -71 845 -37
rect 787 -77 845 -71
rect -887 -142 -841 -118
rect -887 -176 -881 -142
rect -847 -176 -841 -142
rect -887 -214 -841 -176
rect -887 -248 -881 -214
rect -847 -248 -841 -214
rect -887 -286 -841 -248
rect -887 -320 -881 -286
rect -847 -320 -841 -286
rect -887 -358 -841 -320
rect -887 -392 -881 -358
rect -847 -392 -841 -358
rect -887 -430 -841 -392
rect -887 -464 -881 -430
rect -847 -464 -841 -430
rect -887 -502 -841 -464
rect -887 -536 -881 -502
rect -847 -536 -841 -502
rect -887 -560 -841 -536
rect -791 -142 -745 -118
rect -791 -176 -785 -142
rect -751 -176 -745 -142
rect -791 -214 -745 -176
rect -791 -248 -785 -214
rect -751 -248 -745 -214
rect -791 -286 -745 -248
rect -791 -320 -785 -286
rect -751 -320 -745 -286
rect -791 -358 -745 -320
rect -791 -392 -785 -358
rect -751 -392 -745 -358
rect -791 -430 -745 -392
rect -791 -464 -785 -430
rect -751 -464 -745 -430
rect -791 -502 -745 -464
rect -791 -536 -785 -502
rect -751 -536 -745 -502
rect -791 -560 -745 -536
rect -695 -142 -649 -118
rect -695 -176 -689 -142
rect -655 -176 -649 -142
rect -695 -214 -649 -176
rect -695 -248 -689 -214
rect -655 -248 -649 -214
rect -695 -286 -649 -248
rect -695 -320 -689 -286
rect -655 -320 -649 -286
rect -695 -358 -649 -320
rect -695 -392 -689 -358
rect -655 -392 -649 -358
rect -695 -430 -649 -392
rect -695 -464 -689 -430
rect -655 -464 -649 -430
rect -695 -502 -649 -464
rect -695 -536 -689 -502
rect -655 -536 -649 -502
rect -695 -560 -649 -536
rect -599 -142 -553 -118
rect -599 -176 -593 -142
rect -559 -176 -553 -142
rect -599 -214 -553 -176
rect -599 -248 -593 -214
rect -559 -248 -553 -214
rect -599 -286 -553 -248
rect -599 -320 -593 -286
rect -559 -320 -553 -286
rect -599 -358 -553 -320
rect -599 -392 -593 -358
rect -559 -392 -553 -358
rect -599 -430 -553 -392
rect -599 -464 -593 -430
rect -559 -464 -553 -430
rect -599 -502 -553 -464
rect -599 -536 -593 -502
rect -559 -536 -553 -502
rect -599 -560 -553 -536
rect -503 -142 -457 -118
rect -503 -176 -497 -142
rect -463 -176 -457 -142
rect -503 -214 -457 -176
rect -503 -248 -497 -214
rect -463 -248 -457 -214
rect -503 -286 -457 -248
rect -503 -320 -497 -286
rect -463 -320 -457 -286
rect -503 -358 -457 -320
rect -503 -392 -497 -358
rect -463 -392 -457 -358
rect -503 -430 -457 -392
rect -503 -464 -497 -430
rect -463 -464 -457 -430
rect -503 -502 -457 -464
rect -503 -536 -497 -502
rect -463 -536 -457 -502
rect -503 -560 -457 -536
rect -407 -142 -361 -118
rect -407 -176 -401 -142
rect -367 -176 -361 -142
rect -407 -214 -361 -176
rect -407 -248 -401 -214
rect -367 -248 -361 -214
rect -407 -286 -361 -248
rect -407 -320 -401 -286
rect -367 -320 -361 -286
rect -407 -358 -361 -320
rect -407 -392 -401 -358
rect -367 -392 -361 -358
rect -407 -430 -361 -392
rect -407 -464 -401 -430
rect -367 -464 -361 -430
rect -407 -502 -361 -464
rect -407 -536 -401 -502
rect -367 -536 -361 -502
rect -407 -560 -361 -536
rect -311 -142 -265 -118
rect -311 -176 -305 -142
rect -271 -176 -265 -142
rect -311 -214 -265 -176
rect -311 -248 -305 -214
rect -271 -248 -265 -214
rect -311 -286 -265 -248
rect -311 -320 -305 -286
rect -271 -320 -265 -286
rect -311 -358 -265 -320
rect -311 -392 -305 -358
rect -271 -392 -265 -358
rect -311 -430 -265 -392
rect -311 -464 -305 -430
rect -271 -464 -265 -430
rect -311 -502 -265 -464
rect -311 -536 -305 -502
rect -271 -536 -265 -502
rect -311 -560 -265 -536
rect -215 -142 -169 -118
rect -215 -176 -209 -142
rect -175 -176 -169 -142
rect -215 -214 -169 -176
rect -215 -248 -209 -214
rect -175 -248 -169 -214
rect -215 -286 -169 -248
rect -215 -320 -209 -286
rect -175 -320 -169 -286
rect -215 -358 -169 -320
rect -215 -392 -209 -358
rect -175 -392 -169 -358
rect -215 -430 -169 -392
rect -215 -464 -209 -430
rect -175 -464 -169 -430
rect -215 -502 -169 -464
rect -215 -536 -209 -502
rect -175 -536 -169 -502
rect -215 -560 -169 -536
rect -119 -142 -73 -118
rect -119 -176 -113 -142
rect -79 -176 -73 -142
rect -119 -214 -73 -176
rect -119 -248 -113 -214
rect -79 -248 -73 -214
rect -119 -286 -73 -248
rect -119 -320 -113 -286
rect -79 -320 -73 -286
rect -119 -358 -73 -320
rect -119 -392 -113 -358
rect -79 -392 -73 -358
rect -119 -430 -73 -392
rect -119 -464 -113 -430
rect -79 -464 -73 -430
rect -119 -502 -73 -464
rect -119 -536 -113 -502
rect -79 -536 -73 -502
rect -119 -560 -73 -536
rect -23 -142 23 -118
rect -23 -176 -17 -142
rect 17 -176 23 -142
rect -23 -214 23 -176
rect -23 -248 -17 -214
rect 17 -248 23 -214
rect -23 -286 23 -248
rect -23 -320 -17 -286
rect 17 -320 23 -286
rect -23 -358 23 -320
rect -23 -392 -17 -358
rect 17 -392 23 -358
rect -23 -430 23 -392
rect -23 -464 -17 -430
rect 17 -464 23 -430
rect -23 -502 23 -464
rect -23 -536 -17 -502
rect 17 -536 23 -502
rect -23 -560 23 -536
rect 73 -142 119 -118
rect 73 -176 79 -142
rect 113 -176 119 -142
rect 73 -214 119 -176
rect 73 -248 79 -214
rect 113 -248 119 -214
rect 73 -286 119 -248
rect 73 -320 79 -286
rect 113 -320 119 -286
rect 73 -358 119 -320
rect 73 -392 79 -358
rect 113 -392 119 -358
rect 73 -430 119 -392
rect 73 -464 79 -430
rect 113 -464 119 -430
rect 73 -502 119 -464
rect 73 -536 79 -502
rect 113 -536 119 -502
rect 73 -560 119 -536
rect 169 -142 215 -118
rect 169 -176 175 -142
rect 209 -176 215 -142
rect 169 -214 215 -176
rect 169 -248 175 -214
rect 209 -248 215 -214
rect 169 -286 215 -248
rect 169 -320 175 -286
rect 209 -320 215 -286
rect 169 -358 215 -320
rect 169 -392 175 -358
rect 209 -392 215 -358
rect 169 -430 215 -392
rect 169 -464 175 -430
rect 209 -464 215 -430
rect 169 -502 215 -464
rect 169 -536 175 -502
rect 209 -536 215 -502
rect 169 -560 215 -536
rect 265 -142 311 -118
rect 265 -176 271 -142
rect 305 -176 311 -142
rect 265 -214 311 -176
rect 265 -248 271 -214
rect 305 -248 311 -214
rect 265 -286 311 -248
rect 265 -320 271 -286
rect 305 -320 311 -286
rect 265 -358 311 -320
rect 265 -392 271 -358
rect 305 -392 311 -358
rect 265 -430 311 -392
rect 265 -464 271 -430
rect 305 -464 311 -430
rect 265 -502 311 -464
rect 265 -536 271 -502
rect 305 -536 311 -502
rect 265 -560 311 -536
rect 361 -142 407 -118
rect 361 -176 367 -142
rect 401 -176 407 -142
rect 361 -214 407 -176
rect 361 -248 367 -214
rect 401 -248 407 -214
rect 361 -286 407 -248
rect 361 -320 367 -286
rect 401 -320 407 -286
rect 361 -358 407 -320
rect 361 -392 367 -358
rect 401 -392 407 -358
rect 361 -430 407 -392
rect 361 -464 367 -430
rect 401 -464 407 -430
rect 361 -502 407 -464
rect 361 -536 367 -502
rect 401 -536 407 -502
rect 361 -560 407 -536
rect 457 -142 503 -118
rect 457 -176 463 -142
rect 497 -176 503 -142
rect 457 -214 503 -176
rect 457 -248 463 -214
rect 497 -248 503 -214
rect 457 -286 503 -248
rect 457 -320 463 -286
rect 497 -320 503 -286
rect 457 -358 503 -320
rect 457 -392 463 -358
rect 497 -392 503 -358
rect 457 -430 503 -392
rect 457 -464 463 -430
rect 497 -464 503 -430
rect 457 -502 503 -464
rect 457 -536 463 -502
rect 497 -536 503 -502
rect 457 -560 503 -536
rect 553 -142 599 -118
rect 553 -176 559 -142
rect 593 -176 599 -142
rect 553 -214 599 -176
rect 553 -248 559 -214
rect 593 -248 599 -214
rect 553 -286 599 -248
rect 553 -320 559 -286
rect 593 -320 599 -286
rect 553 -358 599 -320
rect 553 -392 559 -358
rect 593 -392 599 -358
rect 553 -430 599 -392
rect 553 -464 559 -430
rect 593 -464 599 -430
rect 553 -502 599 -464
rect 553 -536 559 -502
rect 593 -536 599 -502
rect 553 -560 599 -536
rect 649 -142 695 -118
rect 649 -176 655 -142
rect 689 -176 695 -142
rect 649 -214 695 -176
rect 649 -248 655 -214
rect 689 -248 695 -214
rect 649 -286 695 -248
rect 649 -320 655 -286
rect 689 -320 695 -286
rect 649 -358 695 -320
rect 649 -392 655 -358
rect 689 -392 695 -358
rect 649 -430 695 -392
rect 649 -464 655 -430
rect 689 -464 695 -430
rect 649 -502 695 -464
rect 649 -536 655 -502
rect 689 -536 695 -502
rect 649 -560 695 -536
rect 745 -142 791 -118
rect 745 -176 751 -142
rect 785 -176 791 -142
rect 745 -214 791 -176
rect 745 -248 751 -214
rect 785 -248 791 -214
rect 745 -286 791 -248
rect 745 -320 751 -286
rect 785 -320 791 -286
rect 745 -358 791 -320
rect 745 -392 751 -358
rect 785 -392 791 -358
rect 745 -430 791 -392
rect 745 -464 751 -430
rect 785 -464 791 -430
rect 745 -502 791 -464
rect 745 -536 751 -502
rect 785 -536 791 -502
rect 745 -560 791 -536
rect 841 -142 887 -118
rect 841 -176 847 -142
rect 881 -176 887 -142
rect 841 -214 887 -176
rect 841 -248 847 -214
rect 881 -248 887 -214
rect 841 -286 887 -248
rect 841 -320 847 -286
rect 881 -320 887 -286
rect 841 -358 887 -320
rect 841 -392 847 -358
rect 881 -392 887 -358
rect 841 -430 887 -392
rect 841 -464 847 -430
rect 881 -464 887 -430
rect 841 -502 887 -464
rect 841 -536 847 -502
rect 881 -536 887 -502
rect 841 -560 887 -536
rect -845 -607 -787 -601
rect -845 -641 -833 -607
rect -799 -641 -787 -607
rect -845 -647 -787 -641
rect -653 -607 -595 -601
rect -653 -641 -641 -607
rect -607 -641 -595 -607
rect -653 -647 -595 -641
rect -461 -607 -403 -601
rect -461 -641 -449 -607
rect -415 -641 -403 -607
rect -461 -647 -403 -641
rect -269 -607 -211 -601
rect -269 -641 -257 -607
rect -223 -641 -211 -607
rect -269 -647 -211 -641
rect -77 -607 -19 -601
rect -77 -641 -65 -607
rect -31 -641 -19 -607
rect -77 -647 -19 -641
rect 115 -607 173 -601
rect 115 -641 127 -607
rect 161 -641 173 -607
rect 115 -647 173 -641
rect 307 -607 365 -601
rect 307 -641 319 -607
rect 353 -641 365 -607
rect 307 -647 365 -641
rect 499 -607 557 -601
rect 499 -641 511 -607
rect 545 -641 557 -607
rect 499 -647 557 -641
rect 691 -607 749 -601
rect 691 -641 703 -607
rect 737 -641 749 -607
rect 691 -647 749 -641
<< properties >>
string FIXED_BBOX -978 -726 978 726
<< end >>
