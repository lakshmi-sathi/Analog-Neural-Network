magic
tech sky130A
magscale 1 2
timestamp 1626782926
<< error_p >>
rect -125 681 -67 687
rect 67 681 125 687
rect -125 647 -113 681
rect 67 647 79 681
rect -125 641 -67 647
rect 67 641 125 647
rect -221 -647 -163 -641
rect -29 -647 29 -641
rect 163 -647 221 -641
rect -221 -681 -209 -647
rect -29 -681 -17 -647
rect 163 -681 175 -647
rect -221 -687 -163 -681
rect -29 -687 29 -681
rect 163 -687 221 -681
<< nwell >>
rect -407 -819 407 819
<< pmos >>
rect -207 -600 -177 600
rect -111 -600 -81 600
rect -15 -600 15 600
rect 81 -600 111 600
rect 177 -600 207 600
<< pdiff >>
rect -269 588 -207 600
rect -269 -588 -257 588
rect -223 -588 -207 588
rect -269 -600 -207 -588
rect -177 588 -111 600
rect -177 -588 -161 588
rect -127 -588 -111 588
rect -177 -600 -111 -588
rect -81 588 -15 600
rect -81 -588 -65 588
rect -31 -588 -15 588
rect -81 -600 -15 -588
rect 15 588 81 600
rect 15 -588 31 588
rect 65 -588 81 588
rect 15 -600 81 -588
rect 111 588 177 600
rect 111 -588 127 588
rect 161 -588 177 588
rect 111 -600 177 -588
rect 207 588 269 600
rect 207 -588 223 588
rect 257 -588 269 588
rect 207 -600 269 -588
<< pdiffc >>
rect -257 -588 -223 588
rect -161 -588 -127 588
rect -65 -588 -31 588
rect 31 -588 65 588
rect 127 -588 161 588
rect 223 -588 257 588
<< nsubdiff >>
rect -371 749 -275 783
rect 275 749 371 783
rect -371 687 -337 749
rect 337 687 371 749
rect -371 -749 -337 -687
rect 337 -749 371 -687
rect -371 -783 -275 -749
rect 275 -783 371 -749
<< nsubdiffcont >>
rect -275 749 275 783
rect -371 -687 -337 687
rect 337 -687 371 687
rect -275 -783 275 -749
<< poly >>
rect -129 681 -63 697
rect -129 647 -113 681
rect -79 647 -63 681
rect -129 631 -63 647
rect 63 681 129 697
rect 63 647 79 681
rect 113 647 129 681
rect 63 631 129 647
rect -207 600 -177 626
rect -111 600 -81 631
rect -15 600 15 626
rect 81 600 111 631
rect 177 600 207 626
rect -207 -631 -177 -600
rect -111 -626 -81 -600
rect -15 -631 15 -600
rect 81 -626 111 -600
rect 177 -631 207 -600
rect -225 -647 -159 -631
rect -225 -681 -209 -647
rect -175 -681 -159 -647
rect -225 -697 -159 -681
rect -33 -647 33 -631
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect -33 -697 33 -681
rect 159 -647 225 -631
rect 159 -681 175 -647
rect 209 -681 225 -647
rect 159 -697 225 -681
<< polycont >>
rect -113 647 -79 681
rect 79 647 113 681
rect -209 -681 -175 -647
rect -17 -681 17 -647
rect 175 -681 209 -647
<< locali >>
rect -371 749 -275 783
rect 275 749 371 783
rect -371 687 -337 749
rect 337 687 371 749
rect -129 647 -113 681
rect -79 647 -63 681
rect 63 647 79 681
rect 113 647 129 681
rect -257 588 -223 604
rect -257 -604 -223 -588
rect -161 588 -127 604
rect -161 -604 -127 -588
rect -65 588 -31 604
rect -65 -604 -31 -588
rect 31 588 65 604
rect 31 -604 65 -588
rect 127 588 161 604
rect 127 -604 161 -588
rect 223 588 257 604
rect 223 -604 257 -588
rect -225 -681 -209 -647
rect -175 -681 -159 -647
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect 159 -681 175 -647
rect 209 -681 225 -647
rect -371 -749 -337 -687
rect 337 -749 371 -687
rect -371 -783 -275 -749
rect 275 -783 371 -749
<< viali >>
rect -113 647 -79 681
rect 79 647 113 681
rect -257 -588 -223 588
rect -161 -588 -127 588
rect -65 -588 -31 588
rect 31 -588 65 588
rect 127 -588 161 588
rect 223 -588 257 588
rect -209 -681 -175 -647
rect -17 -681 17 -647
rect 175 -681 209 -647
<< metal1 >>
rect -125 681 -67 687
rect -125 647 -113 681
rect -79 647 -67 681
rect -125 641 -67 647
rect 67 681 125 687
rect 67 647 79 681
rect 113 647 125 681
rect 67 641 125 647
rect -263 588 -217 600
rect -263 -588 -257 588
rect -223 -588 -217 588
rect -263 -600 -217 -588
rect -167 588 -121 600
rect -167 -588 -161 588
rect -127 -588 -121 588
rect -167 -600 -121 -588
rect -71 588 -25 600
rect -71 -588 -65 588
rect -31 -588 -25 588
rect -71 -600 -25 -588
rect 25 588 71 600
rect 25 -588 31 588
rect 65 -588 71 588
rect 25 -600 71 -588
rect 121 588 167 600
rect 121 -588 127 588
rect 161 -588 167 588
rect 121 -600 167 -588
rect 217 588 263 600
rect 217 -588 223 588
rect 257 -588 263 588
rect 217 -600 263 -588
rect -221 -647 -163 -641
rect -221 -681 -209 -647
rect -175 -681 -163 -647
rect -221 -687 -163 -681
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect 17 -681 29 -647
rect -29 -687 29 -681
rect 163 -647 221 -641
rect 163 -681 175 -647
rect 209 -681 221 -647
rect 163 -687 221 -681
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -354 -766 354 766
string parameters w 6 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
