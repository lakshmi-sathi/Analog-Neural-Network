magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 835 35 1267
rect -35 -1267 35 -835
<< xpolyres >>
rect -35 -835 35 835
<< viali >>
rect -17 1213 17 1247
rect -17 1141 17 1175
rect -17 1069 17 1103
rect -17 997 17 1031
rect -17 925 17 959
rect -17 853 17 887
rect -17 -888 17 -854
rect -17 -960 17 -926
rect -17 -1032 17 -998
rect -17 -1104 17 -1070
rect -17 -1176 17 -1142
rect -17 -1248 17 -1214
<< metal1 >>
rect -25 1247 25 1261
rect -25 1213 -17 1247
rect 17 1213 25 1247
rect -25 1175 25 1213
rect -25 1141 -17 1175
rect 17 1141 25 1175
rect -25 1103 25 1141
rect -25 1069 -17 1103
rect 17 1069 25 1103
rect -25 1031 25 1069
rect -25 997 -17 1031
rect 17 997 25 1031
rect -25 959 25 997
rect -25 925 -17 959
rect 17 925 25 959
rect -25 887 25 925
rect -25 853 -17 887
rect 17 853 25 887
rect -25 840 25 853
rect -25 -854 25 -840
rect -25 -888 -17 -854
rect 17 -888 25 -854
rect -25 -926 25 -888
rect -25 -960 -17 -926
rect 17 -960 25 -926
rect -25 -998 25 -960
rect -25 -1032 -17 -998
rect 17 -1032 25 -998
rect -25 -1070 25 -1032
rect -25 -1104 -17 -1070
rect 17 -1104 25 -1070
rect -25 -1142 25 -1104
rect -25 -1176 -17 -1142
rect 17 -1176 25 -1142
rect -25 -1214 25 -1176
rect -25 -1248 -17 -1214
rect 17 -1248 25 -1214
rect -25 -1261 25 -1248
<< end >>
