magic
tech sky130A
magscale 1 2
timestamp 1627838634
<< error_p >>
rect -29 -307 29 -301
rect -29 -341 -17 -307
rect -29 -347 29 -341
<< pwell >>
rect -211 -479 211 479
<< nmos >>
rect -15 -269 15 331
<< ndiff >>
rect -73 319 -15 331
rect -73 -257 -61 319
rect -27 -257 -15 319
rect -73 -269 -15 -257
rect 15 319 73 331
rect 15 -257 27 319
rect 61 -257 73 319
rect 15 -269 73 -257
<< ndiffc >>
rect -61 -257 -27 319
rect 27 -257 61 319
<< psubdiff >>
rect -175 409 -79 443
rect 79 409 175 443
rect -175 347 -141 409
rect 141 347 175 409
rect -175 -409 -141 -347
rect 141 -409 175 -347
rect -175 -443 -79 -409
rect 79 -443 175 -409
<< psubdiffcont >>
rect -79 409 79 443
rect -175 -347 -141 347
rect 141 -347 175 347
rect -79 -443 79 -409
<< poly >>
rect -15 331 15 357
rect -15 -291 15 -269
rect -33 -307 33 -291
rect -33 -341 -17 -307
rect 17 -341 33 -307
rect -33 -357 33 -341
<< polycont >>
rect -17 -341 17 -307
<< locali >>
rect -175 409 -79 443
rect 79 409 175 443
rect -175 347 -141 409
rect 141 347 175 409
rect -61 319 -27 335
rect -61 -273 -27 -257
rect 27 319 61 335
rect 27 -273 61 -257
rect -33 -341 -17 -307
rect 17 -341 33 -307
rect -175 -409 -141 -347
rect 141 -409 175 -347
rect -175 -443 -79 -409
rect 79 -443 175 -409
<< viali >>
rect -61 -257 -27 319
rect 27 -257 61 319
rect -17 -341 17 -307
<< metal1 >>
rect -67 319 -21 331
rect -67 -257 -61 319
rect -27 -257 -21 319
rect -67 -269 -21 -257
rect 21 319 67 331
rect 21 -257 27 319
rect 61 -257 67 319
rect 21 -269 67 -257
rect -29 -307 29 -301
rect -29 -341 -17 -307
rect 17 -341 29 -307
rect -29 -347 29 -341
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -426 158 426
string parameters w 3 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
