magic
tech minimum
magscale 1 2
timestamp 0
<< checkpaint >>
rect 0 0 1 1
<< end >>
