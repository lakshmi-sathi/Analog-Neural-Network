magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 251 35 683
rect -35 -683 35 -251
<< xpolyres >>
rect -35 -251 35 251
<< viali >>
rect -17 629 17 663
rect -17 557 17 591
rect -17 485 17 519
rect -17 413 17 447
rect -17 341 17 375
rect -17 269 17 303
rect -17 -304 17 -270
rect -17 -376 17 -342
rect -17 -448 17 -414
rect -17 -520 17 -486
rect -17 -592 17 -558
rect -17 -664 17 -630
<< metal1 >>
rect -25 663 25 677
rect -25 629 -17 663
rect 17 629 25 663
rect -25 591 25 629
rect -25 557 -17 591
rect 17 557 25 591
rect -25 519 25 557
rect -25 485 -17 519
rect 17 485 25 519
rect -25 447 25 485
rect -25 413 -17 447
rect 17 413 25 447
rect -25 375 25 413
rect -25 341 -17 375
rect 17 341 25 375
rect -25 303 25 341
rect -25 269 -17 303
rect 17 269 25 303
rect -25 256 25 269
rect -25 -270 25 -256
rect -25 -304 -17 -270
rect 17 -304 25 -270
rect -25 -342 25 -304
rect -25 -376 -17 -342
rect 17 -376 25 -342
rect -25 -414 25 -376
rect -25 -448 -17 -414
rect 17 -448 25 -414
rect -25 -486 25 -448
rect -25 -520 -17 -486
rect 17 -520 25 -486
rect -25 -558 25 -520
rect -25 -592 -17 -558
rect 17 -592 25 -558
rect -25 -630 25 -592
rect -25 -664 -17 -630
rect 17 -664 25 -630
rect -25 -677 25 -664
<< end >>
