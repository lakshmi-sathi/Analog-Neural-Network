magic
tech sky130A
magscale 1 2
timestamp 1627115601
<< error_p >>
rect -1901 381 -1843 387
rect -1709 381 -1651 387
rect -1517 381 -1459 387
rect -1325 381 -1267 387
rect -1133 381 -1075 387
rect -941 381 -883 387
rect -749 381 -691 387
rect -557 381 -499 387
rect -365 381 -307 387
rect -173 381 -115 387
rect 19 381 77 387
rect 211 381 269 387
rect 403 381 461 387
rect 595 381 653 387
rect 787 381 845 387
rect 979 381 1037 387
rect 1171 381 1229 387
rect 1363 381 1421 387
rect 1555 381 1613 387
rect 1747 381 1805 387
rect 1939 381 1997 387
rect -1901 347 -1889 381
rect -1709 347 -1697 381
rect -1517 347 -1505 381
rect -1325 347 -1313 381
rect -1133 347 -1121 381
rect -941 347 -929 381
rect -749 347 -737 381
rect -557 347 -545 381
rect -365 347 -353 381
rect -173 347 -161 381
rect 19 347 31 381
rect 211 347 223 381
rect 403 347 415 381
rect 595 347 607 381
rect 787 347 799 381
rect 979 347 991 381
rect 1171 347 1183 381
rect 1363 347 1375 381
rect 1555 347 1567 381
rect 1747 347 1759 381
rect 1939 347 1951 381
rect -1901 341 -1843 347
rect -1709 341 -1651 347
rect -1517 341 -1459 347
rect -1325 341 -1267 347
rect -1133 341 -1075 347
rect -941 341 -883 347
rect -749 341 -691 347
rect -557 341 -499 347
rect -365 341 -307 347
rect -173 341 -115 347
rect 19 341 77 347
rect 211 341 269 347
rect 403 341 461 347
rect 595 341 653 347
rect 787 341 845 347
rect 979 341 1037 347
rect 1171 341 1229 347
rect 1363 341 1421 347
rect 1555 341 1613 347
rect 1747 341 1805 347
rect 1939 341 1997 347
rect -1997 -347 -1939 -341
rect -1805 -347 -1747 -341
rect -1613 -347 -1555 -341
rect -1421 -347 -1363 -341
rect -1229 -347 -1171 -341
rect -1037 -347 -979 -341
rect -845 -347 -787 -341
rect -653 -347 -595 -341
rect -461 -347 -403 -341
rect -269 -347 -211 -341
rect -77 -347 -19 -341
rect 115 -347 173 -341
rect 307 -347 365 -341
rect 499 -347 557 -341
rect 691 -347 749 -341
rect 883 -347 941 -341
rect 1075 -347 1133 -341
rect 1267 -347 1325 -341
rect 1459 -347 1517 -341
rect 1651 -347 1709 -341
rect 1843 -347 1901 -341
rect -1997 -381 -1985 -347
rect -1805 -381 -1793 -347
rect -1613 -381 -1601 -347
rect -1421 -381 -1409 -347
rect -1229 -381 -1217 -347
rect -1037 -381 -1025 -347
rect -845 -381 -833 -347
rect -653 -381 -641 -347
rect -461 -381 -449 -347
rect -269 -381 -257 -347
rect -77 -381 -65 -347
rect 115 -381 127 -347
rect 307 -381 319 -347
rect 499 -381 511 -347
rect 691 -381 703 -347
rect 883 -381 895 -347
rect 1075 -381 1087 -347
rect 1267 -381 1279 -347
rect 1459 -381 1471 -347
rect 1651 -381 1663 -347
rect 1843 -381 1855 -347
rect -1997 -387 -1939 -381
rect -1805 -387 -1747 -381
rect -1613 -387 -1555 -381
rect -1421 -387 -1363 -381
rect -1229 -387 -1171 -381
rect -1037 -387 -979 -381
rect -845 -387 -787 -381
rect -653 -387 -595 -381
rect -461 -387 -403 -381
rect -269 -387 -211 -381
rect -77 -387 -19 -381
rect 115 -387 173 -381
rect 307 -387 365 -381
rect 499 -387 557 -381
rect 691 -387 749 -381
rect 883 -387 941 -381
rect 1075 -387 1133 -381
rect 1267 -387 1325 -381
rect 1459 -387 1517 -381
rect 1651 -387 1709 -381
rect 1843 -387 1901 -381
<< nwell >>
rect -2183 -519 2183 519
<< pmos >>
rect -1983 -300 -1953 300
rect -1887 -300 -1857 300
rect -1791 -300 -1761 300
rect -1695 -300 -1665 300
rect -1599 -300 -1569 300
rect -1503 -300 -1473 300
rect -1407 -300 -1377 300
rect -1311 -300 -1281 300
rect -1215 -300 -1185 300
rect -1119 -300 -1089 300
rect -1023 -300 -993 300
rect -927 -300 -897 300
rect -831 -300 -801 300
rect -735 -300 -705 300
rect -639 -300 -609 300
rect -543 -300 -513 300
rect -447 -300 -417 300
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
rect 417 -300 447 300
rect 513 -300 543 300
rect 609 -300 639 300
rect 705 -300 735 300
rect 801 -300 831 300
rect 897 -300 927 300
rect 993 -300 1023 300
rect 1089 -300 1119 300
rect 1185 -300 1215 300
rect 1281 -300 1311 300
rect 1377 -300 1407 300
rect 1473 -300 1503 300
rect 1569 -300 1599 300
rect 1665 -300 1695 300
rect 1761 -300 1791 300
rect 1857 -300 1887 300
rect 1953 -300 1983 300
<< pdiff >>
rect -2045 288 -1983 300
rect -2045 -288 -2033 288
rect -1999 -288 -1983 288
rect -2045 -300 -1983 -288
rect -1953 288 -1887 300
rect -1953 -288 -1937 288
rect -1903 -288 -1887 288
rect -1953 -300 -1887 -288
rect -1857 288 -1791 300
rect -1857 -288 -1841 288
rect -1807 -288 -1791 288
rect -1857 -300 -1791 -288
rect -1761 288 -1695 300
rect -1761 -288 -1745 288
rect -1711 -288 -1695 288
rect -1761 -300 -1695 -288
rect -1665 288 -1599 300
rect -1665 -288 -1649 288
rect -1615 -288 -1599 288
rect -1665 -300 -1599 -288
rect -1569 288 -1503 300
rect -1569 -288 -1553 288
rect -1519 -288 -1503 288
rect -1569 -300 -1503 -288
rect -1473 288 -1407 300
rect -1473 -288 -1457 288
rect -1423 -288 -1407 288
rect -1473 -300 -1407 -288
rect -1377 288 -1311 300
rect -1377 -288 -1361 288
rect -1327 -288 -1311 288
rect -1377 -300 -1311 -288
rect -1281 288 -1215 300
rect -1281 -288 -1265 288
rect -1231 -288 -1215 288
rect -1281 -300 -1215 -288
rect -1185 288 -1119 300
rect -1185 -288 -1169 288
rect -1135 -288 -1119 288
rect -1185 -300 -1119 -288
rect -1089 288 -1023 300
rect -1089 -288 -1073 288
rect -1039 -288 -1023 288
rect -1089 -300 -1023 -288
rect -993 288 -927 300
rect -993 -288 -977 288
rect -943 -288 -927 288
rect -993 -300 -927 -288
rect -897 288 -831 300
rect -897 -288 -881 288
rect -847 -288 -831 288
rect -897 -300 -831 -288
rect -801 288 -735 300
rect -801 -288 -785 288
rect -751 -288 -735 288
rect -801 -300 -735 -288
rect -705 288 -639 300
rect -705 -288 -689 288
rect -655 -288 -639 288
rect -705 -300 -639 -288
rect -609 288 -543 300
rect -609 -288 -593 288
rect -559 -288 -543 288
rect -609 -300 -543 -288
rect -513 288 -447 300
rect -513 -288 -497 288
rect -463 -288 -447 288
rect -513 -300 -447 -288
rect -417 288 -351 300
rect -417 -288 -401 288
rect -367 -288 -351 288
rect -417 -300 -351 -288
rect -321 288 -255 300
rect -321 -288 -305 288
rect -271 -288 -255 288
rect -321 -300 -255 -288
rect -225 288 -159 300
rect -225 -288 -209 288
rect -175 -288 -159 288
rect -225 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 225 300
rect 159 -288 175 288
rect 209 -288 225 288
rect 159 -300 225 -288
rect 255 288 321 300
rect 255 -288 271 288
rect 305 -288 321 288
rect 255 -300 321 -288
rect 351 288 417 300
rect 351 -288 367 288
rect 401 -288 417 288
rect 351 -300 417 -288
rect 447 288 513 300
rect 447 -288 463 288
rect 497 -288 513 288
rect 447 -300 513 -288
rect 543 288 609 300
rect 543 -288 559 288
rect 593 -288 609 288
rect 543 -300 609 -288
rect 639 288 705 300
rect 639 -288 655 288
rect 689 -288 705 288
rect 639 -300 705 -288
rect 735 288 801 300
rect 735 -288 751 288
rect 785 -288 801 288
rect 735 -300 801 -288
rect 831 288 897 300
rect 831 -288 847 288
rect 881 -288 897 288
rect 831 -300 897 -288
rect 927 288 993 300
rect 927 -288 943 288
rect 977 -288 993 288
rect 927 -300 993 -288
rect 1023 288 1089 300
rect 1023 -288 1039 288
rect 1073 -288 1089 288
rect 1023 -300 1089 -288
rect 1119 288 1185 300
rect 1119 -288 1135 288
rect 1169 -288 1185 288
rect 1119 -300 1185 -288
rect 1215 288 1281 300
rect 1215 -288 1231 288
rect 1265 -288 1281 288
rect 1215 -300 1281 -288
rect 1311 288 1377 300
rect 1311 -288 1327 288
rect 1361 -288 1377 288
rect 1311 -300 1377 -288
rect 1407 288 1473 300
rect 1407 -288 1423 288
rect 1457 -288 1473 288
rect 1407 -300 1473 -288
rect 1503 288 1569 300
rect 1503 -288 1519 288
rect 1553 -288 1569 288
rect 1503 -300 1569 -288
rect 1599 288 1665 300
rect 1599 -288 1615 288
rect 1649 -288 1665 288
rect 1599 -300 1665 -288
rect 1695 288 1761 300
rect 1695 -288 1711 288
rect 1745 -288 1761 288
rect 1695 -300 1761 -288
rect 1791 288 1857 300
rect 1791 -288 1807 288
rect 1841 -288 1857 288
rect 1791 -300 1857 -288
rect 1887 288 1953 300
rect 1887 -288 1903 288
rect 1937 -288 1953 288
rect 1887 -300 1953 -288
rect 1983 288 2045 300
rect 1983 -288 1999 288
rect 2033 -288 2045 288
rect 1983 -300 2045 -288
<< pdiffc >>
rect -2033 -288 -1999 288
rect -1937 -288 -1903 288
rect -1841 -288 -1807 288
rect -1745 -288 -1711 288
rect -1649 -288 -1615 288
rect -1553 -288 -1519 288
rect -1457 -288 -1423 288
rect -1361 -288 -1327 288
rect -1265 -288 -1231 288
rect -1169 -288 -1135 288
rect -1073 -288 -1039 288
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
rect 1039 -288 1073 288
rect 1135 -288 1169 288
rect 1231 -288 1265 288
rect 1327 -288 1361 288
rect 1423 -288 1457 288
rect 1519 -288 1553 288
rect 1615 -288 1649 288
rect 1711 -288 1745 288
rect 1807 -288 1841 288
rect 1903 -288 1937 288
rect 1999 -288 2033 288
<< nsubdiff >>
rect -2147 449 -2051 483
rect 2051 449 2147 483
rect -2147 387 -2113 449
rect 2113 387 2147 449
rect -2147 -449 -2113 -387
rect 2113 -449 2147 -387
rect -2147 -483 -2051 -449
rect 2051 -483 2147 -449
<< nsubdiffcont >>
rect -2051 449 2051 483
rect -2147 -387 -2113 387
rect 2113 -387 2147 387
rect -2051 -483 2051 -449
<< poly >>
rect -1905 381 -1839 397
rect -1905 347 -1889 381
rect -1855 347 -1839 381
rect -1905 331 -1839 347
rect -1713 381 -1647 397
rect -1713 347 -1697 381
rect -1663 347 -1647 381
rect -1713 331 -1647 347
rect -1521 381 -1455 397
rect -1521 347 -1505 381
rect -1471 347 -1455 381
rect -1521 331 -1455 347
rect -1329 381 -1263 397
rect -1329 347 -1313 381
rect -1279 347 -1263 381
rect -1329 331 -1263 347
rect -1137 381 -1071 397
rect -1137 347 -1121 381
rect -1087 347 -1071 381
rect -1137 331 -1071 347
rect -945 381 -879 397
rect -945 347 -929 381
rect -895 347 -879 381
rect -945 331 -879 347
rect -753 381 -687 397
rect -753 347 -737 381
rect -703 347 -687 381
rect -753 331 -687 347
rect -561 381 -495 397
rect -561 347 -545 381
rect -511 347 -495 381
rect -561 331 -495 347
rect -369 381 -303 397
rect -369 347 -353 381
rect -319 347 -303 381
rect -369 331 -303 347
rect -177 381 -111 397
rect -177 347 -161 381
rect -127 347 -111 381
rect -177 331 -111 347
rect 15 381 81 397
rect 15 347 31 381
rect 65 347 81 381
rect 15 331 81 347
rect 207 381 273 397
rect 207 347 223 381
rect 257 347 273 381
rect 207 331 273 347
rect 399 381 465 397
rect 399 347 415 381
rect 449 347 465 381
rect 399 331 465 347
rect 591 381 657 397
rect 591 347 607 381
rect 641 347 657 381
rect 591 331 657 347
rect 783 381 849 397
rect 783 347 799 381
rect 833 347 849 381
rect 783 331 849 347
rect 975 381 1041 397
rect 975 347 991 381
rect 1025 347 1041 381
rect 975 331 1041 347
rect 1167 381 1233 397
rect 1167 347 1183 381
rect 1217 347 1233 381
rect 1167 331 1233 347
rect 1359 381 1425 397
rect 1359 347 1375 381
rect 1409 347 1425 381
rect 1359 331 1425 347
rect 1551 381 1617 397
rect 1551 347 1567 381
rect 1601 347 1617 381
rect 1551 331 1617 347
rect 1743 381 1809 397
rect 1743 347 1759 381
rect 1793 347 1809 381
rect 1743 331 1809 347
rect 1935 381 2001 397
rect 1935 347 1951 381
rect 1985 347 2001 381
rect 1935 331 2001 347
rect -1983 300 -1953 326
rect -1887 300 -1857 331
rect -1791 300 -1761 326
rect -1695 300 -1665 331
rect -1599 300 -1569 326
rect -1503 300 -1473 331
rect -1407 300 -1377 326
rect -1311 300 -1281 331
rect -1215 300 -1185 326
rect -1119 300 -1089 331
rect -1023 300 -993 326
rect -927 300 -897 331
rect -831 300 -801 326
rect -735 300 -705 331
rect -639 300 -609 326
rect -543 300 -513 331
rect -447 300 -417 326
rect -351 300 -321 331
rect -255 300 -225 326
rect -159 300 -129 331
rect -63 300 -33 326
rect 33 300 63 331
rect 129 300 159 326
rect 225 300 255 331
rect 321 300 351 326
rect 417 300 447 331
rect 513 300 543 326
rect 609 300 639 331
rect 705 300 735 326
rect 801 300 831 331
rect 897 300 927 326
rect 993 300 1023 331
rect 1089 300 1119 326
rect 1185 300 1215 331
rect 1281 300 1311 326
rect 1377 300 1407 331
rect 1473 300 1503 326
rect 1569 300 1599 331
rect 1665 300 1695 326
rect 1761 300 1791 331
rect 1857 300 1887 326
rect 1953 300 1983 331
rect -1983 -331 -1953 -300
rect -1887 -326 -1857 -300
rect -1791 -331 -1761 -300
rect -1695 -326 -1665 -300
rect -1599 -331 -1569 -300
rect -1503 -326 -1473 -300
rect -1407 -331 -1377 -300
rect -1311 -326 -1281 -300
rect -1215 -331 -1185 -300
rect -1119 -326 -1089 -300
rect -1023 -331 -993 -300
rect -927 -326 -897 -300
rect -831 -331 -801 -300
rect -735 -326 -705 -300
rect -639 -331 -609 -300
rect -543 -326 -513 -300
rect -447 -331 -417 -300
rect -351 -326 -321 -300
rect -255 -331 -225 -300
rect -159 -326 -129 -300
rect -63 -331 -33 -300
rect 33 -326 63 -300
rect 129 -331 159 -300
rect 225 -326 255 -300
rect 321 -331 351 -300
rect 417 -326 447 -300
rect 513 -331 543 -300
rect 609 -326 639 -300
rect 705 -331 735 -300
rect 801 -326 831 -300
rect 897 -331 927 -300
rect 993 -326 1023 -300
rect 1089 -331 1119 -300
rect 1185 -326 1215 -300
rect 1281 -331 1311 -300
rect 1377 -326 1407 -300
rect 1473 -331 1503 -300
rect 1569 -326 1599 -300
rect 1665 -331 1695 -300
rect 1761 -326 1791 -300
rect 1857 -331 1887 -300
rect 1953 -326 1983 -300
rect -2001 -347 -1935 -331
rect -2001 -381 -1985 -347
rect -1951 -381 -1935 -347
rect -2001 -397 -1935 -381
rect -1809 -347 -1743 -331
rect -1809 -381 -1793 -347
rect -1759 -381 -1743 -347
rect -1809 -397 -1743 -381
rect -1617 -347 -1551 -331
rect -1617 -381 -1601 -347
rect -1567 -381 -1551 -347
rect -1617 -397 -1551 -381
rect -1425 -347 -1359 -331
rect -1425 -381 -1409 -347
rect -1375 -381 -1359 -347
rect -1425 -397 -1359 -381
rect -1233 -347 -1167 -331
rect -1233 -381 -1217 -347
rect -1183 -381 -1167 -347
rect -1233 -397 -1167 -381
rect -1041 -347 -975 -331
rect -1041 -381 -1025 -347
rect -991 -381 -975 -347
rect -1041 -397 -975 -381
rect -849 -347 -783 -331
rect -849 -381 -833 -347
rect -799 -381 -783 -347
rect -849 -397 -783 -381
rect -657 -347 -591 -331
rect -657 -381 -641 -347
rect -607 -381 -591 -347
rect -657 -397 -591 -381
rect -465 -347 -399 -331
rect -465 -381 -449 -347
rect -415 -381 -399 -347
rect -465 -397 -399 -381
rect -273 -347 -207 -331
rect -273 -381 -257 -347
rect -223 -381 -207 -347
rect -273 -397 -207 -381
rect -81 -347 -15 -331
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect -81 -397 -15 -381
rect 111 -347 177 -331
rect 111 -381 127 -347
rect 161 -381 177 -347
rect 111 -397 177 -381
rect 303 -347 369 -331
rect 303 -381 319 -347
rect 353 -381 369 -347
rect 303 -397 369 -381
rect 495 -347 561 -331
rect 495 -381 511 -347
rect 545 -381 561 -347
rect 495 -397 561 -381
rect 687 -347 753 -331
rect 687 -381 703 -347
rect 737 -381 753 -347
rect 687 -397 753 -381
rect 879 -347 945 -331
rect 879 -381 895 -347
rect 929 -381 945 -347
rect 879 -397 945 -381
rect 1071 -347 1137 -331
rect 1071 -381 1087 -347
rect 1121 -381 1137 -347
rect 1071 -397 1137 -381
rect 1263 -347 1329 -331
rect 1263 -381 1279 -347
rect 1313 -381 1329 -347
rect 1263 -397 1329 -381
rect 1455 -347 1521 -331
rect 1455 -381 1471 -347
rect 1505 -381 1521 -347
rect 1455 -397 1521 -381
rect 1647 -347 1713 -331
rect 1647 -381 1663 -347
rect 1697 -381 1713 -347
rect 1647 -397 1713 -381
rect 1839 -347 1905 -331
rect 1839 -381 1855 -347
rect 1889 -381 1905 -347
rect 1839 -397 1905 -381
<< polycont >>
rect -1889 347 -1855 381
rect -1697 347 -1663 381
rect -1505 347 -1471 381
rect -1313 347 -1279 381
rect -1121 347 -1087 381
rect -929 347 -895 381
rect -737 347 -703 381
rect -545 347 -511 381
rect -353 347 -319 381
rect -161 347 -127 381
rect 31 347 65 381
rect 223 347 257 381
rect 415 347 449 381
rect 607 347 641 381
rect 799 347 833 381
rect 991 347 1025 381
rect 1183 347 1217 381
rect 1375 347 1409 381
rect 1567 347 1601 381
rect 1759 347 1793 381
rect 1951 347 1985 381
rect -1985 -381 -1951 -347
rect -1793 -381 -1759 -347
rect -1601 -381 -1567 -347
rect -1409 -381 -1375 -347
rect -1217 -381 -1183 -347
rect -1025 -381 -991 -347
rect -833 -381 -799 -347
rect -641 -381 -607 -347
rect -449 -381 -415 -347
rect -257 -381 -223 -347
rect -65 -381 -31 -347
rect 127 -381 161 -347
rect 319 -381 353 -347
rect 511 -381 545 -347
rect 703 -381 737 -347
rect 895 -381 929 -347
rect 1087 -381 1121 -347
rect 1279 -381 1313 -347
rect 1471 -381 1505 -347
rect 1663 -381 1697 -347
rect 1855 -381 1889 -347
<< locali >>
rect -2147 449 -2051 483
rect 2051 449 2147 483
rect -2147 387 -2113 449
rect 2113 387 2147 449
rect -1905 347 -1889 381
rect -1855 347 -1839 381
rect -1713 347 -1697 381
rect -1663 347 -1647 381
rect -1521 347 -1505 381
rect -1471 347 -1455 381
rect -1329 347 -1313 381
rect -1279 347 -1263 381
rect -1137 347 -1121 381
rect -1087 347 -1071 381
rect -945 347 -929 381
rect -895 347 -879 381
rect -753 347 -737 381
rect -703 347 -687 381
rect -561 347 -545 381
rect -511 347 -495 381
rect -369 347 -353 381
rect -319 347 -303 381
rect -177 347 -161 381
rect -127 347 -111 381
rect 15 347 31 381
rect 65 347 81 381
rect 207 347 223 381
rect 257 347 273 381
rect 399 347 415 381
rect 449 347 465 381
rect 591 347 607 381
rect 641 347 657 381
rect 783 347 799 381
rect 833 347 849 381
rect 975 347 991 381
rect 1025 347 1041 381
rect 1167 347 1183 381
rect 1217 347 1233 381
rect 1359 347 1375 381
rect 1409 347 1425 381
rect 1551 347 1567 381
rect 1601 347 1617 381
rect 1743 347 1759 381
rect 1793 347 1809 381
rect 1935 347 1951 381
rect 1985 347 2001 381
rect -2033 288 -1999 304
rect -2033 -304 -1999 -288
rect -1937 288 -1903 304
rect -1937 -304 -1903 -288
rect -1841 288 -1807 304
rect -1841 -304 -1807 -288
rect -1745 288 -1711 304
rect -1745 -304 -1711 -288
rect -1649 288 -1615 304
rect -1649 -304 -1615 -288
rect -1553 288 -1519 304
rect -1553 -304 -1519 -288
rect -1457 288 -1423 304
rect -1457 -304 -1423 -288
rect -1361 288 -1327 304
rect -1361 -304 -1327 -288
rect -1265 288 -1231 304
rect -1265 -304 -1231 -288
rect -1169 288 -1135 304
rect -1169 -304 -1135 -288
rect -1073 288 -1039 304
rect -1073 -304 -1039 -288
rect -977 288 -943 304
rect -977 -304 -943 -288
rect -881 288 -847 304
rect -881 -304 -847 -288
rect -785 288 -751 304
rect -785 -304 -751 -288
rect -689 288 -655 304
rect -689 -304 -655 -288
rect -593 288 -559 304
rect -593 -304 -559 -288
rect -497 288 -463 304
rect -497 -304 -463 -288
rect -401 288 -367 304
rect -401 -304 -367 -288
rect -305 288 -271 304
rect -305 -304 -271 -288
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect 271 288 305 304
rect 271 -304 305 -288
rect 367 288 401 304
rect 367 -304 401 -288
rect 463 288 497 304
rect 463 -304 497 -288
rect 559 288 593 304
rect 559 -304 593 -288
rect 655 288 689 304
rect 655 -304 689 -288
rect 751 288 785 304
rect 751 -304 785 -288
rect 847 288 881 304
rect 847 -304 881 -288
rect 943 288 977 304
rect 943 -304 977 -288
rect 1039 288 1073 304
rect 1039 -304 1073 -288
rect 1135 288 1169 304
rect 1135 -304 1169 -288
rect 1231 288 1265 304
rect 1231 -304 1265 -288
rect 1327 288 1361 304
rect 1327 -304 1361 -288
rect 1423 288 1457 304
rect 1423 -304 1457 -288
rect 1519 288 1553 304
rect 1519 -304 1553 -288
rect 1615 288 1649 304
rect 1615 -304 1649 -288
rect 1711 288 1745 304
rect 1711 -304 1745 -288
rect 1807 288 1841 304
rect 1807 -304 1841 -288
rect 1903 288 1937 304
rect 1903 -304 1937 -288
rect 1999 288 2033 304
rect 1999 -304 2033 -288
rect -2001 -381 -1985 -347
rect -1951 -381 -1935 -347
rect -1809 -381 -1793 -347
rect -1759 -381 -1743 -347
rect -1617 -381 -1601 -347
rect -1567 -381 -1551 -347
rect -1425 -381 -1409 -347
rect -1375 -381 -1359 -347
rect -1233 -381 -1217 -347
rect -1183 -381 -1167 -347
rect -1041 -381 -1025 -347
rect -991 -381 -975 -347
rect -849 -381 -833 -347
rect -799 -381 -783 -347
rect -657 -381 -641 -347
rect -607 -381 -591 -347
rect -465 -381 -449 -347
rect -415 -381 -399 -347
rect -273 -381 -257 -347
rect -223 -381 -207 -347
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect 111 -381 127 -347
rect 161 -381 177 -347
rect 303 -381 319 -347
rect 353 -381 369 -347
rect 495 -381 511 -347
rect 545 -381 561 -347
rect 687 -381 703 -347
rect 737 -381 753 -347
rect 879 -381 895 -347
rect 929 -381 945 -347
rect 1071 -381 1087 -347
rect 1121 -381 1137 -347
rect 1263 -381 1279 -347
rect 1313 -381 1329 -347
rect 1455 -381 1471 -347
rect 1505 -381 1521 -347
rect 1647 -381 1663 -347
rect 1697 -381 1713 -347
rect 1839 -381 1855 -347
rect 1889 -381 1905 -347
rect -2147 -449 -2113 -387
rect 2113 -449 2147 -387
rect -2147 -483 -2051 -449
rect 2051 -483 2147 -449
<< viali >>
rect -1889 347 -1855 381
rect -1697 347 -1663 381
rect -1505 347 -1471 381
rect -1313 347 -1279 381
rect -1121 347 -1087 381
rect -929 347 -895 381
rect -737 347 -703 381
rect -545 347 -511 381
rect -353 347 -319 381
rect -161 347 -127 381
rect 31 347 65 381
rect 223 347 257 381
rect 415 347 449 381
rect 607 347 641 381
rect 799 347 833 381
rect 991 347 1025 381
rect 1183 347 1217 381
rect 1375 347 1409 381
rect 1567 347 1601 381
rect 1759 347 1793 381
rect 1951 347 1985 381
rect -2033 -288 -1999 288
rect -1937 -288 -1903 288
rect -1841 -288 -1807 288
rect -1745 -288 -1711 288
rect -1649 -288 -1615 288
rect -1553 -288 -1519 288
rect -1457 -288 -1423 288
rect -1361 -288 -1327 288
rect -1265 -288 -1231 288
rect -1169 -288 -1135 288
rect -1073 -288 -1039 288
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
rect 1039 -288 1073 288
rect 1135 -288 1169 288
rect 1231 -288 1265 288
rect 1327 -288 1361 288
rect 1423 -288 1457 288
rect 1519 -288 1553 288
rect 1615 -288 1649 288
rect 1711 -288 1745 288
rect 1807 -288 1841 288
rect 1903 -288 1937 288
rect 1999 -288 2033 288
rect -1985 -381 -1951 -347
rect -1793 -381 -1759 -347
rect -1601 -381 -1567 -347
rect -1409 -381 -1375 -347
rect -1217 -381 -1183 -347
rect -1025 -381 -991 -347
rect -833 -381 -799 -347
rect -641 -381 -607 -347
rect -449 -381 -415 -347
rect -257 -381 -223 -347
rect -65 -381 -31 -347
rect 127 -381 161 -347
rect 319 -381 353 -347
rect 511 -381 545 -347
rect 703 -381 737 -347
rect 895 -381 929 -347
rect 1087 -381 1121 -347
rect 1279 -381 1313 -347
rect 1471 -381 1505 -347
rect 1663 -381 1697 -347
rect 1855 -381 1889 -347
<< metal1 >>
rect -1901 381 -1843 387
rect -1901 347 -1889 381
rect -1855 347 -1843 381
rect -1901 341 -1843 347
rect -1709 381 -1651 387
rect -1709 347 -1697 381
rect -1663 347 -1651 381
rect -1709 341 -1651 347
rect -1517 381 -1459 387
rect -1517 347 -1505 381
rect -1471 347 -1459 381
rect -1517 341 -1459 347
rect -1325 381 -1267 387
rect -1325 347 -1313 381
rect -1279 347 -1267 381
rect -1325 341 -1267 347
rect -1133 381 -1075 387
rect -1133 347 -1121 381
rect -1087 347 -1075 381
rect -1133 341 -1075 347
rect -941 381 -883 387
rect -941 347 -929 381
rect -895 347 -883 381
rect -941 341 -883 347
rect -749 381 -691 387
rect -749 347 -737 381
rect -703 347 -691 381
rect -749 341 -691 347
rect -557 381 -499 387
rect -557 347 -545 381
rect -511 347 -499 381
rect -557 341 -499 347
rect -365 381 -307 387
rect -365 347 -353 381
rect -319 347 -307 381
rect -365 341 -307 347
rect -173 381 -115 387
rect -173 347 -161 381
rect -127 347 -115 381
rect -173 341 -115 347
rect 19 381 77 387
rect 19 347 31 381
rect 65 347 77 381
rect 19 341 77 347
rect 211 381 269 387
rect 211 347 223 381
rect 257 347 269 381
rect 211 341 269 347
rect 403 381 461 387
rect 403 347 415 381
rect 449 347 461 381
rect 403 341 461 347
rect 595 381 653 387
rect 595 347 607 381
rect 641 347 653 381
rect 595 341 653 347
rect 787 381 845 387
rect 787 347 799 381
rect 833 347 845 381
rect 787 341 845 347
rect 979 381 1037 387
rect 979 347 991 381
rect 1025 347 1037 381
rect 979 341 1037 347
rect 1171 381 1229 387
rect 1171 347 1183 381
rect 1217 347 1229 381
rect 1171 341 1229 347
rect 1363 381 1421 387
rect 1363 347 1375 381
rect 1409 347 1421 381
rect 1363 341 1421 347
rect 1555 381 1613 387
rect 1555 347 1567 381
rect 1601 347 1613 381
rect 1555 341 1613 347
rect 1747 381 1805 387
rect 1747 347 1759 381
rect 1793 347 1805 381
rect 1747 341 1805 347
rect 1939 381 1997 387
rect 1939 347 1951 381
rect 1985 347 1997 381
rect 1939 341 1997 347
rect -2039 288 -1993 300
rect -2039 -288 -2033 288
rect -1999 -288 -1993 288
rect -2039 -300 -1993 -288
rect -1943 288 -1897 300
rect -1943 -288 -1937 288
rect -1903 -288 -1897 288
rect -1943 -300 -1897 -288
rect -1847 288 -1801 300
rect -1847 -288 -1841 288
rect -1807 -288 -1801 288
rect -1847 -300 -1801 -288
rect -1751 288 -1705 300
rect -1751 -288 -1745 288
rect -1711 -288 -1705 288
rect -1751 -300 -1705 -288
rect -1655 288 -1609 300
rect -1655 -288 -1649 288
rect -1615 -288 -1609 288
rect -1655 -300 -1609 -288
rect -1559 288 -1513 300
rect -1559 -288 -1553 288
rect -1519 -288 -1513 288
rect -1559 -300 -1513 -288
rect -1463 288 -1417 300
rect -1463 -288 -1457 288
rect -1423 -288 -1417 288
rect -1463 -300 -1417 -288
rect -1367 288 -1321 300
rect -1367 -288 -1361 288
rect -1327 -288 -1321 288
rect -1367 -300 -1321 -288
rect -1271 288 -1225 300
rect -1271 -288 -1265 288
rect -1231 -288 -1225 288
rect -1271 -300 -1225 -288
rect -1175 288 -1129 300
rect -1175 -288 -1169 288
rect -1135 -288 -1129 288
rect -1175 -300 -1129 -288
rect -1079 288 -1033 300
rect -1079 -288 -1073 288
rect -1039 -288 -1033 288
rect -1079 -300 -1033 -288
rect -983 288 -937 300
rect -983 -288 -977 288
rect -943 -288 -937 288
rect -983 -300 -937 -288
rect -887 288 -841 300
rect -887 -288 -881 288
rect -847 -288 -841 288
rect -887 -300 -841 -288
rect -791 288 -745 300
rect -791 -288 -785 288
rect -751 -288 -745 288
rect -791 -300 -745 -288
rect -695 288 -649 300
rect -695 -288 -689 288
rect -655 -288 -649 288
rect -695 -300 -649 -288
rect -599 288 -553 300
rect -599 -288 -593 288
rect -559 -288 -553 288
rect -599 -300 -553 -288
rect -503 288 -457 300
rect -503 -288 -497 288
rect -463 -288 -457 288
rect -503 -300 -457 -288
rect -407 288 -361 300
rect -407 -288 -401 288
rect -367 -288 -361 288
rect -407 -300 -361 -288
rect -311 288 -265 300
rect -311 -288 -305 288
rect -271 -288 -265 288
rect -311 -300 -265 -288
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect 265 288 311 300
rect 265 -288 271 288
rect 305 -288 311 288
rect 265 -300 311 -288
rect 361 288 407 300
rect 361 -288 367 288
rect 401 -288 407 288
rect 361 -300 407 -288
rect 457 288 503 300
rect 457 -288 463 288
rect 497 -288 503 288
rect 457 -300 503 -288
rect 553 288 599 300
rect 553 -288 559 288
rect 593 -288 599 288
rect 553 -300 599 -288
rect 649 288 695 300
rect 649 -288 655 288
rect 689 -288 695 288
rect 649 -300 695 -288
rect 745 288 791 300
rect 745 -288 751 288
rect 785 -288 791 288
rect 745 -300 791 -288
rect 841 288 887 300
rect 841 -288 847 288
rect 881 -288 887 288
rect 841 -300 887 -288
rect 937 288 983 300
rect 937 -288 943 288
rect 977 -288 983 288
rect 937 -300 983 -288
rect 1033 288 1079 300
rect 1033 -288 1039 288
rect 1073 -288 1079 288
rect 1033 -300 1079 -288
rect 1129 288 1175 300
rect 1129 -288 1135 288
rect 1169 -288 1175 288
rect 1129 -300 1175 -288
rect 1225 288 1271 300
rect 1225 -288 1231 288
rect 1265 -288 1271 288
rect 1225 -300 1271 -288
rect 1321 288 1367 300
rect 1321 -288 1327 288
rect 1361 -288 1367 288
rect 1321 -300 1367 -288
rect 1417 288 1463 300
rect 1417 -288 1423 288
rect 1457 -288 1463 288
rect 1417 -300 1463 -288
rect 1513 288 1559 300
rect 1513 -288 1519 288
rect 1553 -288 1559 288
rect 1513 -300 1559 -288
rect 1609 288 1655 300
rect 1609 -288 1615 288
rect 1649 -288 1655 288
rect 1609 -300 1655 -288
rect 1705 288 1751 300
rect 1705 -288 1711 288
rect 1745 -288 1751 288
rect 1705 -300 1751 -288
rect 1801 288 1847 300
rect 1801 -288 1807 288
rect 1841 -288 1847 288
rect 1801 -300 1847 -288
rect 1897 288 1943 300
rect 1897 -288 1903 288
rect 1937 -288 1943 288
rect 1897 -300 1943 -288
rect 1993 288 2039 300
rect 1993 -288 1999 288
rect 2033 -288 2039 288
rect 1993 -300 2039 -288
rect -1997 -347 -1939 -341
rect -1997 -381 -1985 -347
rect -1951 -381 -1939 -347
rect -1997 -387 -1939 -381
rect -1805 -347 -1747 -341
rect -1805 -381 -1793 -347
rect -1759 -381 -1747 -347
rect -1805 -387 -1747 -381
rect -1613 -347 -1555 -341
rect -1613 -381 -1601 -347
rect -1567 -381 -1555 -347
rect -1613 -387 -1555 -381
rect -1421 -347 -1363 -341
rect -1421 -381 -1409 -347
rect -1375 -381 -1363 -347
rect -1421 -387 -1363 -381
rect -1229 -347 -1171 -341
rect -1229 -381 -1217 -347
rect -1183 -381 -1171 -347
rect -1229 -387 -1171 -381
rect -1037 -347 -979 -341
rect -1037 -381 -1025 -347
rect -991 -381 -979 -347
rect -1037 -387 -979 -381
rect -845 -347 -787 -341
rect -845 -381 -833 -347
rect -799 -381 -787 -347
rect -845 -387 -787 -381
rect -653 -347 -595 -341
rect -653 -381 -641 -347
rect -607 -381 -595 -347
rect -653 -387 -595 -381
rect -461 -347 -403 -341
rect -461 -381 -449 -347
rect -415 -381 -403 -347
rect -461 -387 -403 -381
rect -269 -347 -211 -341
rect -269 -381 -257 -347
rect -223 -381 -211 -347
rect -269 -387 -211 -381
rect -77 -347 -19 -341
rect -77 -381 -65 -347
rect -31 -381 -19 -347
rect -77 -387 -19 -381
rect 115 -347 173 -341
rect 115 -381 127 -347
rect 161 -381 173 -347
rect 115 -387 173 -381
rect 307 -347 365 -341
rect 307 -381 319 -347
rect 353 -381 365 -347
rect 307 -387 365 -381
rect 499 -347 557 -341
rect 499 -381 511 -347
rect 545 -381 557 -347
rect 499 -387 557 -381
rect 691 -347 749 -341
rect 691 -381 703 -347
rect 737 -381 749 -347
rect 691 -387 749 -381
rect 883 -347 941 -341
rect 883 -381 895 -347
rect 929 -381 941 -347
rect 883 -387 941 -381
rect 1075 -347 1133 -341
rect 1075 -381 1087 -347
rect 1121 -381 1133 -347
rect 1075 -387 1133 -381
rect 1267 -347 1325 -341
rect 1267 -381 1279 -347
rect 1313 -381 1325 -347
rect 1267 -387 1325 -381
rect 1459 -347 1517 -341
rect 1459 -381 1471 -347
rect 1505 -381 1517 -347
rect 1459 -387 1517 -381
rect 1651 -347 1709 -341
rect 1651 -381 1663 -347
rect 1697 -381 1709 -347
rect 1651 -387 1709 -381
rect 1843 -347 1901 -341
rect 1843 -381 1855 -347
rect 1889 -381 1901 -347
rect 1843 -387 1901 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -2130 -466 2130 466
string parameters w 3 l 0.15 m 1 nf 42 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
