magic
tech sky130A
magscale 1 2
timestamp 1627836603
<< pwell >>
rect 10446 320 10450 334
<< locali >>
rect 2558 1138 2565 1160
rect 2479 1125 2513 1129
rect 2527 1125 2561 1131
rect 2479 1012 2561 1125
rect 2190 978 2561 1012
rect 8149 200 8369 234
rect 8165 173 8369 200
rect 8335 102 8369 173
rect 8334 18 8530 102
<< viali >>
rect 126 726 224 1630
<< metal1 >>
rect 2316 2400 2960 2430
rect 2316 2374 3294 2400
rect 134 1650 236 1654
rect 108 1632 236 1650
rect 108 1630 270 1632
rect 108 1108 126 1630
rect -1354 382 -932 776
rect -762 726 126 1108
rect 224 1108 270 1630
rect 2316 1450 2456 2374
rect 2816 2352 3294 2374
rect 2816 2350 2958 2352
rect 2250 1432 2456 1450
rect 2250 1132 2272 1432
rect 2386 1270 2456 1432
rect 3956 1378 4044 1384
rect 4246 1378 4300 1992
rect 4429 1378 4483 1989
rect 4623 1378 4677 1981
rect 4823 1378 4877 1969
rect 5011 1378 5065 1969
rect 5207 1378 5261 1963
rect 5387 1378 5441 1985
rect 5583 1378 5637 1963
rect 5779 1378 5833 1965
rect 5975 1378 6029 1967
rect 6155 1378 6209 1969
rect 6355 1378 6409 1969
rect 6551 1378 6605 1977
rect 6739 1378 6793 1973
rect 7754 1491 7948 1492
rect 8260 1491 8443 1493
rect 7754 1474 8443 1491
rect 7390 1453 8443 1474
rect 7390 1426 7948 1453
rect 2386 1182 2498 1270
rect 3956 1242 3968 1378
rect 6824 1242 6834 1378
rect 3956 1236 4094 1242
rect 2386 1132 2412 1182
rect 2250 1114 2412 1132
rect 224 726 352 1108
rect 4042 744 4094 1236
rect 4234 744 4286 1242
rect 4430 744 4482 1242
rect 4614 744 4666 1242
rect 4806 744 4858 1242
rect 5004 744 5056 1242
rect 5196 744 5248 1242
rect 5388 744 5440 1242
rect 5580 744 5632 1242
rect 5776 744 5828 1242
rect 5964 744 6016 1242
rect 6160 744 6212 1242
rect 6344 744 6396 1242
rect 8260 936 8443 1453
rect 8260 898 8444 936
rect -762 710 352 726
rect -306 706 210 710
rect 8260 582 8290 898
rect 8422 582 8444 898
rect 10412 686 10656 1630
rect -1346 -46 -924 118
rect -762 60 -340 454
rect 8260 400 8444 582
rect 8258 344 8444 400
rect 8224 256 8444 344
rect -10 234 0 238
rect -194 -46 0 234
rect 156 -46 166 238
rect -1346 -54 78 -46
rect -1346 -142 -32 -54
<< via1 >>
rect 2272 1132 2386 1432
rect 3968 1242 6824 1378
rect 8290 582 8422 898
rect 0 -46 156 238
<< metal2 >>
rect 66 2780 10696 2910
rect 254 2666 2318 2780
rect 2455 2560 4030 2680
rect 2455 2559 3822 2560
rect 3880 1947 4030 2560
rect 3880 1797 4032 1947
rect 3881 1760 4032 1797
rect 4156 1760 8268 1762
rect 3881 1742 8268 1760
rect 3881 1626 4108 1742
rect 8208 1626 8268 1742
rect 3881 1612 8268 1626
rect 3881 1611 4143 1612
rect 3881 1609 4031 1611
rect 2258 1432 2400 1444
rect 2258 1430 2272 1432
rect 2386 1430 2400 1432
rect 2258 1132 2270 1430
rect 2390 1132 2400 1430
rect 3962 1378 6824 1388
rect 3962 1242 3968 1378
rect 3962 1232 6824 1242
rect 2258 1120 2400 1132
rect 3708 1054 3812 1084
rect 4006 1054 6848 1064
rect 3708 1048 6848 1054
rect 3708 932 4006 1048
rect 6650 932 6848 1048
rect 3708 926 6848 932
rect 4006 918 6848 926
rect 0 238 156 248
rect 6701 197 6847 918
rect 8276 898 8434 906
rect 8276 582 8290 898
rect 8422 582 8434 898
rect 8276 570 8434 582
rect 6701 146 6850 197
rect 6701 141 6868 146
rect 6701 51 8240 141
rect 6702 -5 8240 51
rect 6702 -8 6888 -5
rect 0 -56 156 -46
rect 94 -234 10724 -104
<< via2 >>
rect 4108 1626 8208 1742
rect 2270 1132 2272 1430
rect 2272 1132 2386 1430
rect 2386 1132 2390 1430
rect 3968 1242 6824 1378
rect 4006 932 6650 1048
rect 0 -46 156 238
rect 8292 594 8414 888
<< metal3 >>
rect 4162 1760 8274 1846
rect 4068 1742 8274 1760
rect 4068 1626 4108 1742
rect 8208 1688 8274 1742
rect 8208 1626 8264 1688
rect 4068 1608 8264 1626
rect 2182 1430 2400 1480
rect 2182 1132 2270 1430
rect 2390 1132 2400 1430
rect 3902 1383 4044 1384
rect 3902 1378 6834 1383
rect 3902 1362 3968 1378
rect 3708 1266 3968 1362
rect 3902 1242 3968 1266
rect 6824 1242 6834 1378
rect 3902 1237 6834 1242
rect 3902 1236 4044 1237
rect 2182 1102 2400 1132
rect 4006 1056 6672 1064
rect 4000 1048 6672 1056
rect 4000 932 4006 1048
rect 6650 932 6672 1048
rect 4000 918 6672 932
rect 8272 1052 8580 1148
rect 4000 880 6448 918
rect 4004 860 6448 880
rect 8272 888 8590 1052
rect 8272 594 8292 888
rect 8414 594 8436 888
rect 8272 556 8436 594
rect -10 238 166 243
rect -10 -46 0 238
rect 156 -46 166 238
rect 10518 232 10702 262
rect 6926 194 7020 198
rect 6918 44 6928 194
rect 7020 44 7030 194
rect 6926 40 7020 44
rect -10 -51 166 -46
rect 10518 -30 10540 232
rect 10668 -30 10702 232
rect 10518 -72 10702 -30
<< via3 >>
rect 0 -46 156 238
rect 6928 44 7020 194
rect 10540 -30 10668 232
<< metal4 >>
rect -15 238 10686 244
rect -15 -46 0 238
rect 156 232 10686 238
rect 156 194 10540 232
rect 156 44 6928 194
rect 7020 44 10540 194
rect 156 -30 10540 44
rect 10668 -30 10686 232
rect 156 -46 10686 -30
rect -15 -54 10686 -46
use biaspmos  biaspmos_0
timestamp 1627800606
transform 1 0 4116 0 1 3370
box -52 -1706 4314 -516
use Stage2_inv  Stage2_inv_0
timestamp 1627803151
transform 1 0 2512 0 1 1150
box -102 -170 1308 1530
use Stage2_inv  Stage2_inv_1
timestamp 1627803151
transform -1 0 8210 0 1 224
box -102 -170 1308 1530
use biasnmos  biasnmos_0
timestamp 1627800883
transform 1 0 2416 0 1 90
box -106 -320 4260 833
use Stage1_inv  Stage1_inv_1
timestamp 1627668659
transform -1 0 10370 0 1 1184
box -166 -1292 1986 1598
use Stage1_inv  Stage1_inv_0
timestamp 1627668659
transform 1 0 362 0 1 1178
box -166 -1292 1986 1598
use sky130_fd_pr__res_xhigh_po_0p35_NZHUVC  sky130_fd_pr__res_xhigh_po_0p35_NZHUVC_0
timestamp 1627748178
transform 0 1 -842 -1 0 741
box -37 -508 37 508
use sky130_fd_pr__res_xhigh_po_0p35_NZHUVC  sky130_fd_pr__res_xhigh_po_0p35_NZHUVC_1
timestamp 1627748178
transform 0 1 -844 -1 0 423
box -37 -508 37 508
use sky130_fd_pr__res_xhigh_po_0p35_NZHUVC  sky130_fd_pr__res_xhigh_po_0p35_NZHUVC_2
timestamp 1627748178
transform 0 1 -840 -1 0 93
box -37 -508 37 508
<< labels >>
rlabel metal1 10448 716 10622 1604 1 in2
port 4 n
rlabel metal2 110 -220 10712 -114 1 GND
port 2 n
rlabel metal2 78 2790 10680 2896 1 VDD
port 1 n
rlabel metal1 126 728 222 1632 1 in1
port 6 n
rlabel metal1 -748 722 100 1096 1 in
port 7 n
rlabel metal3 10526 -62 10694 254 1 out
port 8 n
<< end >>
