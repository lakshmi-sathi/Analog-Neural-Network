magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_p >>
rect -29 83 29 89
rect -29 49 -17 83
rect -29 43 29 49
<< nmos >>
rect -15 -73 15 11
<< ndiff >>
rect -73 -14 -15 11
rect -73 -48 -61 -14
rect -27 -48 -15 -14
rect -73 -73 -15 -48
rect 15 -14 73 11
rect 15 -48 27 -14
rect 61 -48 73 -14
rect 15 -73 73 -48
<< ndiffc >>
rect -61 -48 -27 -14
rect 27 -48 61 -14
<< poly >>
rect -33 83 33 99
rect -33 49 -17 83
rect 17 49 33 83
rect -33 33 33 49
rect -15 11 15 33
rect -15 -99 15 -73
<< polycont >>
rect -17 49 17 83
<< locali >>
rect -33 49 -17 83
rect 17 49 33 83
rect -61 -14 -27 15
rect -61 -77 -27 -48
rect 27 -14 61 15
rect 27 -77 61 -48
<< viali >>
rect -17 49 17 83
rect -61 -48 -27 -14
rect 27 -48 61 -14
<< metal1 >>
rect -29 83 29 89
rect -29 49 -17 83
rect 17 49 29 83
rect -29 43 29 49
rect -67 -14 -21 11
rect -67 -48 -61 -14
rect -27 -48 -21 -14
rect -67 -73 -21 -48
rect 21 -14 67 11
rect 21 -48 27 -14
rect 61 -48 67 -14
rect 21 -73 67 -48
<< end >>
