magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< nwell >>
rect -24 -640 4314 -636
rect -52 -1438 4314 -640
rect -52 -1442 348 -1438
<< pwell >>
rect 252 -1706 2310 -1502
<< psubdiff >>
rect 252 -1519 2310 -1502
rect 252 -1689 278 -1519
rect 2284 -1689 2310 -1519
rect 252 -1706 2310 -1689
<< nsubdiff >>
rect -16 -713 32 -682
rect -16 -747 -10 -713
rect 24 -747 32 -713
rect -16 -781 32 -747
rect -16 -815 -10 -781
rect 24 -815 32 -781
rect -16 -849 32 -815
rect -16 -883 -10 -849
rect 24 -883 32 -849
rect -16 -917 32 -883
rect -16 -951 -10 -917
rect 24 -951 32 -917
rect -16 -985 32 -951
rect -16 -1019 -10 -985
rect 24 -1019 32 -985
rect -16 -1053 32 -1019
rect -16 -1087 -10 -1053
rect 24 -1087 32 -1053
rect -16 -1121 32 -1087
rect -16 -1155 -10 -1121
rect 24 -1155 32 -1121
rect -16 -1189 32 -1155
rect -16 -1223 -10 -1189
rect 24 -1223 32 -1189
rect -16 -1257 32 -1223
rect -16 -1291 -10 -1257
rect 24 -1291 32 -1257
rect -16 -1325 32 -1291
rect -16 -1359 -10 -1325
rect 24 -1359 32 -1325
rect 4230 -709 4278 -678
rect 4230 -743 4236 -709
rect 4270 -743 4278 -709
rect 4230 -777 4278 -743
rect 4230 -811 4236 -777
rect 4270 -811 4278 -777
rect 4230 -845 4278 -811
rect 4230 -879 4236 -845
rect 4270 -879 4278 -845
rect 4230 -913 4278 -879
rect 4230 -947 4236 -913
rect 4270 -947 4278 -913
rect 4230 -981 4278 -947
rect 4230 -1015 4236 -981
rect 4270 -1015 4278 -981
rect 4230 -1049 4278 -1015
rect 4230 -1083 4236 -1049
rect 4270 -1083 4278 -1049
rect 4230 -1117 4278 -1083
rect 4230 -1151 4236 -1117
rect 4270 -1151 4278 -1117
rect 4230 -1185 4278 -1151
rect 4230 -1219 4236 -1185
rect 4270 -1219 4278 -1185
rect 4230 -1253 4278 -1219
rect 4230 -1287 4236 -1253
rect 4270 -1287 4278 -1253
rect 4230 -1321 4278 -1287
rect -16 -1390 32 -1359
rect 4230 -1355 4236 -1321
rect 4270 -1355 4278 -1321
rect 4230 -1386 4278 -1355
<< psubdiffcont >>
rect 278 -1689 2284 -1519
<< nsubdiffcont >>
rect -10 -747 24 -713
rect -10 -815 24 -781
rect -10 -883 24 -849
rect -10 -951 24 -917
rect -10 -1019 24 -985
rect -10 -1087 24 -1053
rect -10 -1155 24 -1121
rect -10 -1223 24 -1189
rect -10 -1291 24 -1257
rect -10 -1359 24 -1325
rect 4236 -743 4270 -709
rect 4236 -811 4270 -777
rect 4236 -879 4270 -845
rect 4236 -947 4270 -913
rect 4236 -1015 4270 -981
rect 4236 -1083 4270 -1049
rect 4236 -1151 4270 -1117
rect 4236 -1219 4270 -1185
rect 4236 -1287 4270 -1253
rect 4236 -1355 4270 -1321
<< poly >>
rect 4084 -1393 4114 -1341
rect 4027 -1423 4114 -1393
<< locali >>
rect 88 -551 4166 -538
rect 88 -585 131 -551
rect 165 -585 203 -551
rect 237 -585 275 -551
rect 309 -585 347 -551
rect 381 -585 419 -551
rect 453 -585 491 -551
rect 525 -585 563 -551
rect 597 -585 635 -551
rect 669 -585 707 -551
rect 741 -585 779 -551
rect 813 -585 851 -551
rect 885 -585 923 -551
rect 957 -585 995 -551
rect 1029 -585 1067 -551
rect 1101 -585 1139 -551
rect 1173 -585 1211 -551
rect 1245 -585 1283 -551
rect 1317 -585 1355 -551
rect 1389 -585 1427 -551
rect 1461 -585 1499 -551
rect 1533 -585 1571 -551
rect 1605 -585 1643 -551
rect 1677 -585 1715 -551
rect 1749 -585 1787 -551
rect 1821 -585 1859 -551
rect 1893 -585 1931 -551
rect 1965 -585 2003 -551
rect 2037 -585 2075 -551
rect 2109 -585 2147 -551
rect 2181 -585 2219 -551
rect 2253 -585 2291 -551
rect 2325 -585 2363 -551
rect 2397 -585 2435 -551
rect 2469 -585 2507 -551
rect 2541 -585 2579 -551
rect 2613 -585 2651 -551
rect 2685 -585 2723 -551
rect 2757 -585 2795 -551
rect 2829 -585 2867 -551
rect 2901 -585 2939 -551
rect 2973 -585 3011 -551
rect 3045 -585 3083 -551
rect 3117 -585 3155 -551
rect 3189 -585 3227 -551
rect 3261 -585 3299 -551
rect 3333 -585 3371 -551
rect 3405 -585 3443 -551
rect 3477 -585 3515 -551
rect 3549 -585 3587 -551
rect 3621 -585 3659 -551
rect 3693 -585 3731 -551
rect 3765 -585 3803 -551
rect 3837 -585 3875 -551
rect 3909 -585 3947 -551
rect 3981 -585 4019 -551
rect 4053 -585 4091 -551
rect 4125 -585 4166 -551
rect 88 -600 4166 -585
rect -16 -713 32 -682
rect -16 -747 -10 -713
rect 24 -747 32 -713
rect -16 -781 32 -747
rect -16 -815 -10 -781
rect 24 -815 32 -781
rect -16 -849 32 -815
rect -16 -883 -10 -849
rect 24 -883 32 -849
rect -16 -917 32 -883
rect -16 -951 -10 -917
rect 24 -951 32 -917
rect -16 -985 32 -951
rect -16 -1019 -10 -985
rect 24 -1019 32 -985
rect -16 -1053 32 -1019
rect -16 -1087 -10 -1053
rect 24 -1087 32 -1053
rect -16 -1121 32 -1087
rect -16 -1155 -10 -1121
rect 24 -1155 32 -1121
rect -16 -1189 32 -1155
rect -16 -1223 -10 -1189
rect 24 -1223 32 -1189
rect -16 -1257 32 -1223
rect -16 -1291 -10 -1257
rect 24 -1291 32 -1257
rect -16 -1325 32 -1291
rect -16 -1359 -10 -1325
rect 24 -1359 32 -1325
rect -16 -1390 32 -1359
rect 4230 -709 4278 -678
rect 4230 -743 4236 -709
rect 4270 -743 4278 -709
rect 4230 -777 4278 -743
rect 4230 -811 4236 -777
rect 4270 -811 4278 -777
rect 4230 -845 4278 -811
rect 4230 -879 4236 -845
rect 4270 -879 4278 -845
rect 4230 -913 4278 -879
rect 4230 -947 4236 -913
rect 4270 -947 4278 -913
rect 4230 -981 4278 -947
rect 4230 -1015 4236 -981
rect 4270 -1015 4278 -981
rect 4230 -1049 4278 -1015
rect 4230 -1083 4236 -1049
rect 4270 -1083 4278 -1049
rect 4230 -1117 4278 -1083
rect 4230 -1151 4236 -1117
rect 4270 -1151 4278 -1117
rect 4230 -1185 4278 -1151
rect 4230 -1219 4236 -1185
rect 4270 -1219 4278 -1185
rect 4230 -1253 4278 -1219
rect 4230 -1287 4236 -1253
rect 4270 -1287 4278 -1253
rect 4230 -1321 4278 -1287
rect 4230 -1355 4236 -1321
rect 4270 -1355 4278 -1321
rect 4230 -1386 4278 -1355
rect 260 -1519 2302 -1502
rect 260 -1689 278 -1519
rect 2284 -1689 2302 -1519
rect 260 -1706 2302 -1689
<< viali >>
rect 131 -585 165 -551
rect 203 -585 237 -551
rect 275 -585 309 -551
rect 347 -585 381 -551
rect 419 -585 453 -551
rect 491 -585 525 -551
rect 563 -585 597 -551
rect 635 -585 669 -551
rect 707 -585 741 -551
rect 779 -585 813 -551
rect 851 -585 885 -551
rect 923 -585 957 -551
rect 995 -585 1029 -551
rect 1067 -585 1101 -551
rect 1139 -585 1173 -551
rect 1211 -585 1245 -551
rect 1283 -585 1317 -551
rect 1355 -585 1389 -551
rect 1427 -585 1461 -551
rect 1499 -585 1533 -551
rect 1571 -585 1605 -551
rect 1643 -585 1677 -551
rect 1715 -585 1749 -551
rect 1787 -585 1821 -551
rect 1859 -585 1893 -551
rect 1931 -585 1965 -551
rect 2003 -585 2037 -551
rect 2075 -585 2109 -551
rect 2147 -585 2181 -551
rect 2219 -585 2253 -551
rect 2291 -585 2325 -551
rect 2363 -585 2397 -551
rect 2435 -585 2469 -551
rect 2507 -585 2541 -551
rect 2579 -585 2613 -551
rect 2651 -585 2685 -551
rect 2723 -585 2757 -551
rect 2795 -585 2829 -551
rect 2867 -585 2901 -551
rect 2939 -585 2973 -551
rect 3011 -585 3045 -551
rect 3083 -585 3117 -551
rect 3155 -585 3189 -551
rect 3227 -585 3261 -551
rect 3299 -585 3333 -551
rect 3371 -585 3405 -551
rect 3443 -585 3477 -551
rect 3515 -585 3549 -551
rect 3587 -585 3621 -551
rect 3659 -585 3693 -551
rect 3731 -585 3765 -551
rect 3803 -585 3837 -551
rect 3875 -585 3909 -551
rect 3947 -585 3981 -551
rect 4019 -585 4053 -551
rect 4091 -585 4125 -551
<< metal1 >>
rect 84 -540 4172 -538
rect 84 -592 118 -540
rect 170 -592 182 -540
rect 234 -551 246 -540
rect 298 -551 310 -540
rect 362 -551 374 -540
rect 426 -551 438 -540
rect 490 -551 502 -540
rect 554 -551 566 -540
rect 237 -585 246 -551
rect 309 -585 310 -551
rect 490 -585 491 -551
rect 554 -585 563 -551
rect 234 -592 246 -585
rect 298 -592 310 -585
rect 362 -592 374 -585
rect 426 -592 438 -585
rect 490 -592 502 -585
rect 554 -592 566 -585
rect 618 -592 630 -540
rect 682 -592 694 -540
rect 746 -592 758 -540
rect 810 -551 822 -540
rect 874 -551 886 -540
rect 938 -551 950 -540
rect 1002 -551 1014 -540
rect 1066 -551 1078 -540
rect 1130 -551 1142 -540
rect 813 -585 822 -551
rect 885 -585 886 -551
rect 1066 -585 1067 -551
rect 1130 -585 1139 -551
rect 810 -592 822 -585
rect 874 -592 886 -585
rect 938 -592 950 -585
rect 1002 -592 1014 -585
rect 1066 -592 1078 -585
rect 1130 -592 1142 -585
rect 1194 -592 1206 -540
rect 1258 -592 1270 -540
rect 1322 -592 1334 -540
rect 1386 -551 1398 -540
rect 1450 -551 1462 -540
rect 1514 -551 1526 -540
rect 1578 -551 1590 -540
rect 1642 -551 1654 -540
rect 1706 -551 1718 -540
rect 1389 -585 1398 -551
rect 1461 -585 1462 -551
rect 1642 -585 1643 -551
rect 1706 -585 1715 -551
rect 1386 -592 1398 -585
rect 1450 -592 1462 -585
rect 1514 -592 1526 -585
rect 1578 -592 1590 -585
rect 1642 -592 1654 -585
rect 1706 -592 1718 -585
rect 1770 -592 1782 -540
rect 1834 -592 1846 -540
rect 1898 -592 1910 -540
rect 1962 -551 1974 -540
rect 2026 -551 2038 -540
rect 2090 -551 2102 -540
rect 2154 -551 2166 -540
rect 2218 -551 2230 -540
rect 2282 -551 2294 -540
rect 1965 -585 1974 -551
rect 2037 -585 2038 -551
rect 2218 -585 2219 -551
rect 2282 -585 2291 -551
rect 1962 -592 1974 -585
rect 2026 -592 2038 -585
rect 2090 -592 2102 -585
rect 2154 -592 2166 -585
rect 2218 -592 2230 -585
rect 2282 -592 2294 -585
rect 2346 -592 2358 -540
rect 2410 -592 2422 -540
rect 2474 -592 2486 -540
rect 2538 -551 2550 -540
rect 2602 -551 2614 -540
rect 2666 -551 2678 -540
rect 2730 -551 2742 -540
rect 2794 -551 2806 -540
rect 2858 -551 2870 -540
rect 2541 -585 2550 -551
rect 2613 -585 2614 -551
rect 2794 -585 2795 -551
rect 2858 -585 2867 -551
rect 2538 -592 2550 -585
rect 2602 -592 2614 -585
rect 2666 -592 2678 -585
rect 2730 -592 2742 -585
rect 2794 -592 2806 -585
rect 2858 -592 2870 -585
rect 2922 -592 2934 -540
rect 2986 -592 2998 -540
rect 3050 -592 3062 -540
rect 3114 -551 3126 -540
rect 3178 -551 3190 -540
rect 3242 -551 3254 -540
rect 3306 -551 3318 -540
rect 3370 -551 3382 -540
rect 3434 -551 3446 -540
rect 3117 -585 3126 -551
rect 3189 -585 3190 -551
rect 3370 -585 3371 -551
rect 3434 -585 3443 -551
rect 3114 -592 3126 -585
rect 3178 -592 3190 -585
rect 3242 -592 3254 -585
rect 3306 -592 3318 -585
rect 3370 -592 3382 -585
rect 3434 -592 3446 -585
rect 3498 -592 3510 -540
rect 3562 -592 3574 -540
rect 3626 -592 3638 -540
rect 3690 -551 3702 -540
rect 3754 -551 3766 -540
rect 3818 -551 3830 -540
rect 3882 -551 3894 -540
rect 3946 -551 3958 -540
rect 4010 -551 4022 -540
rect 3693 -585 3702 -551
rect 3765 -585 3766 -551
rect 3946 -585 3947 -551
rect 4010 -585 4019 -551
rect 3690 -592 3702 -585
rect 3754 -592 3766 -585
rect 3818 -592 3830 -585
rect 3882 -592 3894 -585
rect 3946 -592 3958 -585
rect 4010 -592 4022 -585
rect 4074 -592 4086 -540
rect 4138 -592 4172 -540
rect 84 -604 4172 -592
rect 226 -650 4130 -642
rect 226 -704 4132 -650
rect 226 -706 4130 -704
rect 82 -765 150 -742
rect 82 -817 90 -765
rect 142 -817 150 -765
rect 82 -829 150 -817
rect 82 -881 90 -829
rect 142 -881 150 -829
rect 82 -893 150 -881
rect 82 -945 90 -893
rect 142 -945 150 -893
rect 82 -957 150 -945
rect 82 -1009 90 -957
rect 142 -1009 150 -957
rect 82 -1032 150 -1009
rect 274 -765 342 -742
rect 274 -817 282 -765
rect 334 -817 342 -765
rect 274 -829 342 -817
rect 274 -881 282 -829
rect 334 -881 342 -829
rect 274 -893 342 -881
rect 274 -945 282 -893
rect 334 -945 342 -893
rect 274 -957 342 -945
rect 274 -1009 282 -957
rect 334 -1009 342 -957
rect 274 -1032 342 -1009
rect 466 -765 534 -742
rect 466 -817 474 -765
rect 526 -817 534 -765
rect 466 -829 534 -817
rect 466 -881 474 -829
rect 526 -881 534 -829
rect 466 -893 534 -881
rect 466 -945 474 -893
rect 526 -945 534 -893
rect 466 -957 534 -945
rect 466 -1009 474 -957
rect 526 -1009 534 -957
rect 466 -1032 534 -1009
rect 658 -765 726 -742
rect 658 -817 666 -765
rect 718 -817 726 -765
rect 658 -829 726 -817
rect 658 -881 666 -829
rect 718 -881 726 -829
rect 658 -893 726 -881
rect 658 -945 666 -893
rect 718 -945 726 -893
rect 658 -957 726 -945
rect 658 -1009 666 -957
rect 718 -1009 726 -957
rect 658 -1032 726 -1009
rect 850 -765 918 -742
rect 850 -817 858 -765
rect 910 -817 918 -765
rect 850 -829 918 -817
rect 850 -881 858 -829
rect 910 -881 918 -829
rect 850 -893 918 -881
rect 850 -945 858 -893
rect 910 -945 918 -893
rect 850 -957 918 -945
rect 850 -1009 858 -957
rect 910 -1009 918 -957
rect 850 -1032 918 -1009
rect 1042 -765 1110 -742
rect 1042 -817 1050 -765
rect 1102 -817 1110 -765
rect 1042 -829 1110 -817
rect 1042 -881 1050 -829
rect 1102 -881 1110 -829
rect 1042 -893 1110 -881
rect 1042 -945 1050 -893
rect 1102 -945 1110 -893
rect 1042 -957 1110 -945
rect 1042 -1009 1050 -957
rect 1102 -1009 1110 -957
rect 1042 -1032 1110 -1009
rect 1234 -765 1302 -742
rect 1234 -817 1242 -765
rect 1294 -817 1302 -765
rect 1234 -829 1302 -817
rect 1234 -881 1242 -829
rect 1294 -881 1302 -829
rect 1234 -893 1302 -881
rect 1234 -945 1242 -893
rect 1294 -945 1302 -893
rect 1234 -957 1302 -945
rect 1234 -1009 1242 -957
rect 1294 -1009 1302 -957
rect 1234 -1032 1302 -1009
rect 1426 -765 1494 -742
rect 1426 -817 1434 -765
rect 1486 -817 1494 -765
rect 1426 -829 1494 -817
rect 1426 -881 1434 -829
rect 1486 -881 1494 -829
rect 1426 -893 1494 -881
rect 1426 -945 1434 -893
rect 1486 -945 1494 -893
rect 1426 -957 1494 -945
rect 1426 -1009 1434 -957
rect 1486 -1009 1494 -957
rect 1426 -1032 1494 -1009
rect 1618 -765 1686 -742
rect 1618 -817 1626 -765
rect 1678 -817 1686 -765
rect 1618 -829 1686 -817
rect 1618 -881 1626 -829
rect 1678 -881 1686 -829
rect 1618 -893 1686 -881
rect 1618 -945 1626 -893
rect 1678 -945 1686 -893
rect 1618 -957 1686 -945
rect 1618 -1009 1626 -957
rect 1678 -1009 1686 -957
rect 1618 -1032 1686 -1009
rect 1810 -765 1878 -742
rect 1810 -817 1818 -765
rect 1870 -817 1878 -765
rect 1810 -829 1878 -817
rect 1810 -881 1818 -829
rect 1870 -881 1878 -829
rect 1810 -893 1878 -881
rect 1810 -945 1818 -893
rect 1870 -945 1878 -893
rect 1810 -957 1878 -945
rect 1810 -1009 1818 -957
rect 1870 -1009 1878 -957
rect 1810 -1032 1878 -1009
rect 2002 -765 2070 -742
rect 2002 -817 2010 -765
rect 2062 -817 2070 -765
rect 2002 -829 2070 -817
rect 2002 -881 2010 -829
rect 2062 -881 2070 -829
rect 2002 -893 2070 -881
rect 2002 -945 2010 -893
rect 2062 -945 2070 -893
rect 2002 -957 2070 -945
rect 2002 -1009 2010 -957
rect 2062 -1009 2070 -957
rect 2002 -1032 2070 -1009
rect 2194 -765 2262 -742
rect 2194 -817 2202 -765
rect 2254 -817 2262 -765
rect 2194 -829 2262 -817
rect 2194 -881 2202 -829
rect 2254 -881 2262 -829
rect 2194 -893 2262 -881
rect 2194 -945 2202 -893
rect 2254 -945 2262 -893
rect 2194 -957 2262 -945
rect 2194 -1009 2202 -957
rect 2254 -1009 2262 -957
rect 2194 -1032 2262 -1009
rect 2386 -765 2454 -742
rect 2386 -817 2394 -765
rect 2446 -817 2454 -765
rect 2386 -829 2454 -817
rect 2386 -881 2394 -829
rect 2446 -881 2454 -829
rect 2386 -893 2454 -881
rect 2386 -945 2394 -893
rect 2446 -945 2454 -893
rect 2386 -957 2454 -945
rect 2386 -1009 2394 -957
rect 2446 -1009 2454 -957
rect 2386 -1032 2454 -1009
rect 2578 -765 2646 -742
rect 2578 -817 2586 -765
rect 2638 -817 2646 -765
rect 2578 -829 2646 -817
rect 2578 -881 2586 -829
rect 2638 -881 2646 -829
rect 2578 -893 2646 -881
rect 2578 -945 2586 -893
rect 2638 -945 2646 -893
rect 2578 -957 2646 -945
rect 2578 -1009 2586 -957
rect 2638 -1009 2646 -957
rect 2578 -1032 2646 -1009
rect 2770 -765 2838 -742
rect 2770 -817 2778 -765
rect 2830 -817 2838 -765
rect 2770 -829 2838 -817
rect 2770 -881 2778 -829
rect 2830 -881 2838 -829
rect 2770 -893 2838 -881
rect 2770 -945 2778 -893
rect 2830 -945 2838 -893
rect 2770 -957 2838 -945
rect 2770 -1009 2778 -957
rect 2830 -1009 2838 -957
rect 2770 -1032 2838 -1009
rect 2962 -765 3030 -742
rect 2962 -817 2970 -765
rect 3022 -817 3030 -765
rect 2962 -829 3030 -817
rect 2962 -881 2970 -829
rect 3022 -881 3030 -829
rect 2962 -893 3030 -881
rect 2962 -945 2970 -893
rect 3022 -945 3030 -893
rect 2962 -957 3030 -945
rect 2962 -1009 2970 -957
rect 3022 -1009 3030 -957
rect 2962 -1032 3030 -1009
rect 3154 -765 3222 -742
rect 3154 -817 3162 -765
rect 3214 -817 3222 -765
rect 3154 -829 3222 -817
rect 3154 -881 3162 -829
rect 3214 -881 3222 -829
rect 3154 -893 3222 -881
rect 3154 -945 3162 -893
rect 3214 -945 3222 -893
rect 3154 -957 3222 -945
rect 3154 -1009 3162 -957
rect 3214 -1009 3222 -957
rect 3154 -1032 3222 -1009
rect 3346 -765 3414 -742
rect 3346 -817 3354 -765
rect 3406 -817 3414 -765
rect 3346 -829 3414 -817
rect 3346 -881 3354 -829
rect 3406 -881 3414 -829
rect 3346 -893 3414 -881
rect 3346 -945 3354 -893
rect 3406 -945 3414 -893
rect 3346 -957 3414 -945
rect 3346 -1009 3354 -957
rect 3406 -1009 3414 -957
rect 3346 -1032 3414 -1009
rect 3538 -765 3606 -742
rect 3538 -817 3546 -765
rect 3598 -817 3606 -765
rect 3538 -829 3606 -817
rect 3538 -881 3546 -829
rect 3598 -881 3606 -829
rect 3538 -893 3606 -881
rect 3538 -945 3546 -893
rect 3598 -945 3606 -893
rect 3538 -957 3606 -945
rect 3538 -1009 3546 -957
rect 3598 -1009 3606 -957
rect 3538 -1032 3606 -1009
rect 3730 -765 3798 -742
rect 3730 -817 3738 -765
rect 3790 -817 3798 -765
rect 3730 -829 3798 -817
rect 3730 -881 3738 -829
rect 3790 -881 3798 -829
rect 3730 -893 3798 -881
rect 3730 -945 3738 -893
rect 3790 -945 3798 -893
rect 3730 -957 3798 -945
rect 3730 -1009 3738 -957
rect 3790 -1009 3798 -957
rect 3730 -1032 3798 -1009
rect 3922 -765 3990 -742
rect 3922 -817 3930 -765
rect 3982 -817 3990 -765
rect 3922 -829 3990 -817
rect 3922 -881 3930 -829
rect 3982 -881 3990 -829
rect 3922 -893 3990 -881
rect 3922 -945 3930 -893
rect 3982 -945 3990 -893
rect 3922 -957 3990 -945
rect 3922 -1009 3930 -957
rect 3982 -1009 3990 -957
rect 3922 -1032 3990 -1009
rect 4114 -765 4182 -742
rect 4114 -817 4122 -765
rect 4174 -817 4182 -765
rect 4114 -829 4182 -817
rect 4114 -881 4122 -829
rect 4174 -881 4182 -829
rect 4114 -893 4182 -881
rect 4114 -945 4122 -893
rect 4174 -945 4182 -893
rect 4114 -957 4182 -945
rect 4114 -1009 4122 -957
rect 4174 -1009 4182 -957
rect 4114 -1032 4182 -1009
rect 180 -1089 244 -1080
rect 180 -1141 186 -1089
rect 238 -1141 244 -1089
rect 180 -1153 244 -1141
rect 180 -1205 186 -1153
rect 238 -1205 244 -1153
rect 180 -1217 244 -1205
rect 180 -1269 186 -1217
rect 238 -1269 244 -1217
rect 180 -1281 244 -1269
rect 180 -1333 186 -1281
rect 238 -1333 244 -1281
rect 180 -1350 244 -1333
rect 372 -1089 436 -1080
rect 372 -1141 378 -1089
rect 430 -1141 436 -1089
rect 372 -1153 436 -1141
rect 372 -1205 378 -1153
rect 430 -1205 436 -1153
rect 372 -1217 436 -1205
rect 372 -1269 378 -1217
rect 430 -1269 436 -1217
rect 372 -1281 436 -1269
rect 372 -1333 378 -1281
rect 430 -1333 436 -1281
rect 372 -1350 436 -1333
rect 564 -1089 628 -1080
rect 564 -1141 570 -1089
rect 622 -1141 628 -1089
rect 564 -1153 628 -1141
rect 564 -1205 570 -1153
rect 622 -1205 628 -1153
rect 564 -1217 628 -1205
rect 564 -1269 570 -1217
rect 622 -1269 628 -1217
rect 564 -1281 628 -1269
rect 564 -1333 570 -1281
rect 622 -1333 628 -1281
rect 564 -1350 628 -1333
rect 756 -1089 820 -1080
rect 756 -1141 762 -1089
rect 814 -1141 820 -1089
rect 756 -1153 820 -1141
rect 756 -1205 762 -1153
rect 814 -1205 820 -1153
rect 756 -1217 820 -1205
rect 756 -1269 762 -1217
rect 814 -1269 820 -1217
rect 756 -1281 820 -1269
rect 756 -1333 762 -1281
rect 814 -1333 820 -1281
rect 756 -1350 820 -1333
rect 948 -1089 1012 -1080
rect 948 -1141 954 -1089
rect 1006 -1141 1012 -1089
rect 948 -1153 1012 -1141
rect 948 -1205 954 -1153
rect 1006 -1205 1012 -1153
rect 948 -1217 1012 -1205
rect 948 -1269 954 -1217
rect 1006 -1269 1012 -1217
rect 948 -1281 1012 -1269
rect 948 -1333 954 -1281
rect 1006 -1333 1012 -1281
rect 948 -1350 1012 -1333
rect 1140 -1089 1204 -1080
rect 1140 -1141 1146 -1089
rect 1198 -1141 1204 -1089
rect 1140 -1153 1204 -1141
rect 1140 -1205 1146 -1153
rect 1198 -1205 1204 -1153
rect 1140 -1217 1204 -1205
rect 1140 -1269 1146 -1217
rect 1198 -1269 1204 -1217
rect 1140 -1281 1204 -1269
rect 1140 -1333 1146 -1281
rect 1198 -1333 1204 -1281
rect 1140 -1350 1204 -1333
rect 1332 -1089 1396 -1080
rect 1332 -1141 1338 -1089
rect 1390 -1141 1396 -1089
rect 1332 -1153 1396 -1141
rect 1332 -1205 1338 -1153
rect 1390 -1205 1396 -1153
rect 1332 -1217 1396 -1205
rect 1332 -1269 1338 -1217
rect 1390 -1269 1396 -1217
rect 1332 -1281 1396 -1269
rect 1332 -1333 1338 -1281
rect 1390 -1333 1396 -1281
rect 1332 -1350 1396 -1333
rect 1524 -1089 1588 -1080
rect 1524 -1141 1530 -1089
rect 1582 -1141 1588 -1089
rect 1524 -1153 1588 -1141
rect 1524 -1205 1530 -1153
rect 1582 -1205 1588 -1153
rect 1524 -1217 1588 -1205
rect 1524 -1269 1530 -1217
rect 1582 -1269 1588 -1217
rect 1524 -1281 1588 -1269
rect 1524 -1333 1530 -1281
rect 1582 -1333 1588 -1281
rect 1524 -1350 1588 -1333
rect 1716 -1089 1780 -1080
rect 1716 -1141 1722 -1089
rect 1774 -1141 1780 -1089
rect 1716 -1153 1780 -1141
rect 1716 -1205 1722 -1153
rect 1774 -1205 1780 -1153
rect 1716 -1217 1780 -1205
rect 1716 -1269 1722 -1217
rect 1774 -1269 1780 -1217
rect 1716 -1281 1780 -1269
rect 1716 -1333 1722 -1281
rect 1774 -1333 1780 -1281
rect 1716 -1350 1780 -1333
rect 1908 -1089 1972 -1080
rect 1908 -1141 1914 -1089
rect 1966 -1141 1972 -1089
rect 1908 -1153 1972 -1141
rect 1908 -1205 1914 -1153
rect 1966 -1205 1972 -1153
rect 1908 -1217 1972 -1205
rect 1908 -1269 1914 -1217
rect 1966 -1269 1972 -1217
rect 1908 -1281 1972 -1269
rect 1908 -1333 1914 -1281
rect 1966 -1333 1972 -1281
rect 1908 -1350 1972 -1333
rect 2100 -1089 2164 -1080
rect 2100 -1141 2106 -1089
rect 2158 -1141 2164 -1089
rect 2100 -1153 2164 -1141
rect 2100 -1205 2106 -1153
rect 2158 -1205 2164 -1153
rect 2100 -1217 2164 -1205
rect 2100 -1269 2106 -1217
rect 2158 -1269 2164 -1217
rect 2100 -1281 2164 -1269
rect 2100 -1333 2106 -1281
rect 2158 -1333 2164 -1281
rect 2100 -1350 2164 -1333
rect 2292 -1089 2356 -1080
rect 2292 -1141 2298 -1089
rect 2350 -1141 2356 -1089
rect 2292 -1153 2356 -1141
rect 2292 -1205 2298 -1153
rect 2350 -1205 2356 -1153
rect 2292 -1217 2356 -1205
rect 2292 -1269 2298 -1217
rect 2350 -1269 2356 -1217
rect 2292 -1281 2356 -1269
rect 2292 -1333 2298 -1281
rect 2350 -1333 2356 -1281
rect 2292 -1350 2356 -1333
rect 2484 -1089 2548 -1080
rect 2484 -1141 2490 -1089
rect 2542 -1141 2548 -1089
rect 2484 -1153 2548 -1141
rect 2484 -1205 2490 -1153
rect 2542 -1205 2548 -1153
rect 2484 -1217 2548 -1205
rect 2484 -1269 2490 -1217
rect 2542 -1269 2548 -1217
rect 2484 -1281 2548 -1269
rect 2484 -1333 2490 -1281
rect 2542 -1333 2548 -1281
rect 2484 -1350 2548 -1333
rect 2676 -1089 2740 -1080
rect 2676 -1141 2682 -1089
rect 2734 -1141 2740 -1089
rect 2676 -1153 2740 -1141
rect 2676 -1205 2682 -1153
rect 2734 -1205 2740 -1153
rect 2676 -1217 2740 -1205
rect 2676 -1269 2682 -1217
rect 2734 -1269 2740 -1217
rect 2676 -1281 2740 -1269
rect 2676 -1333 2682 -1281
rect 2734 -1333 2740 -1281
rect 2676 -1350 2740 -1333
rect 2868 -1089 2932 -1080
rect 2868 -1141 2874 -1089
rect 2926 -1141 2932 -1089
rect 2868 -1153 2932 -1141
rect 2868 -1205 2874 -1153
rect 2926 -1205 2932 -1153
rect 2868 -1217 2932 -1205
rect 2868 -1269 2874 -1217
rect 2926 -1269 2932 -1217
rect 2868 -1281 2932 -1269
rect 2868 -1333 2874 -1281
rect 2926 -1333 2932 -1281
rect 2868 -1350 2932 -1333
rect 3060 -1089 3124 -1080
rect 3060 -1141 3066 -1089
rect 3118 -1141 3124 -1089
rect 3060 -1153 3124 -1141
rect 3060 -1205 3066 -1153
rect 3118 -1205 3124 -1153
rect 3060 -1217 3124 -1205
rect 3060 -1269 3066 -1217
rect 3118 -1269 3124 -1217
rect 3060 -1281 3124 -1269
rect 3060 -1333 3066 -1281
rect 3118 -1333 3124 -1281
rect 3060 -1350 3124 -1333
rect 3252 -1089 3316 -1080
rect 3252 -1141 3258 -1089
rect 3310 -1141 3316 -1089
rect 3252 -1153 3316 -1141
rect 3252 -1205 3258 -1153
rect 3310 -1205 3316 -1153
rect 3252 -1217 3316 -1205
rect 3252 -1269 3258 -1217
rect 3310 -1269 3316 -1217
rect 3252 -1281 3316 -1269
rect 3252 -1333 3258 -1281
rect 3310 -1333 3316 -1281
rect 3252 -1350 3316 -1333
rect 3444 -1089 3508 -1080
rect 3444 -1141 3450 -1089
rect 3502 -1141 3508 -1089
rect 3444 -1153 3508 -1141
rect 3444 -1205 3450 -1153
rect 3502 -1205 3508 -1153
rect 3444 -1217 3508 -1205
rect 3444 -1269 3450 -1217
rect 3502 -1269 3508 -1217
rect 3444 -1281 3508 -1269
rect 3444 -1333 3450 -1281
rect 3502 -1333 3508 -1281
rect 3444 -1350 3508 -1333
rect 3636 -1089 3700 -1080
rect 3636 -1141 3642 -1089
rect 3694 -1141 3700 -1089
rect 3636 -1153 3700 -1141
rect 3636 -1205 3642 -1153
rect 3694 -1205 3700 -1153
rect 3636 -1217 3700 -1205
rect 3636 -1269 3642 -1217
rect 3694 -1269 3700 -1217
rect 3636 -1281 3700 -1269
rect 3636 -1333 3642 -1281
rect 3694 -1333 3700 -1281
rect 3636 -1350 3700 -1333
rect 3828 -1089 3892 -1080
rect 3828 -1141 3834 -1089
rect 3886 -1141 3892 -1089
rect 3828 -1153 3892 -1141
rect 3828 -1205 3834 -1153
rect 3886 -1205 3892 -1153
rect 3828 -1217 3892 -1205
rect 3828 -1269 3834 -1217
rect 3886 -1269 3892 -1217
rect 3828 -1281 3892 -1269
rect 3828 -1333 3834 -1281
rect 3886 -1333 3892 -1281
rect 3828 -1350 3892 -1333
rect 4020 -1089 4084 -1080
rect 4020 -1141 4026 -1089
rect 4078 -1141 4084 -1089
rect 4020 -1153 4084 -1141
rect 4020 -1205 4026 -1153
rect 4078 -1205 4084 -1153
rect 4020 -1217 4084 -1205
rect 4020 -1269 4026 -1217
rect 4078 -1269 4084 -1217
rect 4020 -1281 4084 -1269
rect 4020 -1333 4026 -1281
rect 4078 -1333 4084 -1281
rect 4020 -1350 4084 -1333
rect 132 -1432 4036 -1378
<< via1 >>
rect 118 -551 170 -540
rect 118 -585 131 -551
rect 131 -585 165 -551
rect 165 -585 170 -551
rect 118 -592 170 -585
rect 182 -551 234 -540
rect 246 -551 298 -540
rect 310 -551 362 -540
rect 374 -551 426 -540
rect 438 -551 490 -540
rect 502 -551 554 -540
rect 566 -551 618 -540
rect 182 -585 203 -551
rect 203 -585 234 -551
rect 246 -585 275 -551
rect 275 -585 298 -551
rect 310 -585 347 -551
rect 347 -585 362 -551
rect 374 -585 381 -551
rect 381 -585 419 -551
rect 419 -585 426 -551
rect 438 -585 453 -551
rect 453 -585 490 -551
rect 502 -585 525 -551
rect 525 -585 554 -551
rect 566 -585 597 -551
rect 597 -585 618 -551
rect 182 -592 234 -585
rect 246 -592 298 -585
rect 310 -592 362 -585
rect 374 -592 426 -585
rect 438 -592 490 -585
rect 502 -592 554 -585
rect 566 -592 618 -585
rect 630 -551 682 -540
rect 630 -585 635 -551
rect 635 -585 669 -551
rect 669 -585 682 -551
rect 630 -592 682 -585
rect 694 -551 746 -540
rect 694 -585 707 -551
rect 707 -585 741 -551
rect 741 -585 746 -551
rect 694 -592 746 -585
rect 758 -551 810 -540
rect 822 -551 874 -540
rect 886 -551 938 -540
rect 950 -551 1002 -540
rect 1014 -551 1066 -540
rect 1078 -551 1130 -540
rect 1142 -551 1194 -540
rect 758 -585 779 -551
rect 779 -585 810 -551
rect 822 -585 851 -551
rect 851 -585 874 -551
rect 886 -585 923 -551
rect 923 -585 938 -551
rect 950 -585 957 -551
rect 957 -585 995 -551
rect 995 -585 1002 -551
rect 1014 -585 1029 -551
rect 1029 -585 1066 -551
rect 1078 -585 1101 -551
rect 1101 -585 1130 -551
rect 1142 -585 1173 -551
rect 1173 -585 1194 -551
rect 758 -592 810 -585
rect 822 -592 874 -585
rect 886 -592 938 -585
rect 950 -592 1002 -585
rect 1014 -592 1066 -585
rect 1078 -592 1130 -585
rect 1142 -592 1194 -585
rect 1206 -551 1258 -540
rect 1206 -585 1211 -551
rect 1211 -585 1245 -551
rect 1245 -585 1258 -551
rect 1206 -592 1258 -585
rect 1270 -551 1322 -540
rect 1270 -585 1283 -551
rect 1283 -585 1317 -551
rect 1317 -585 1322 -551
rect 1270 -592 1322 -585
rect 1334 -551 1386 -540
rect 1398 -551 1450 -540
rect 1462 -551 1514 -540
rect 1526 -551 1578 -540
rect 1590 -551 1642 -540
rect 1654 -551 1706 -540
rect 1718 -551 1770 -540
rect 1334 -585 1355 -551
rect 1355 -585 1386 -551
rect 1398 -585 1427 -551
rect 1427 -585 1450 -551
rect 1462 -585 1499 -551
rect 1499 -585 1514 -551
rect 1526 -585 1533 -551
rect 1533 -585 1571 -551
rect 1571 -585 1578 -551
rect 1590 -585 1605 -551
rect 1605 -585 1642 -551
rect 1654 -585 1677 -551
rect 1677 -585 1706 -551
rect 1718 -585 1749 -551
rect 1749 -585 1770 -551
rect 1334 -592 1386 -585
rect 1398 -592 1450 -585
rect 1462 -592 1514 -585
rect 1526 -592 1578 -585
rect 1590 -592 1642 -585
rect 1654 -592 1706 -585
rect 1718 -592 1770 -585
rect 1782 -551 1834 -540
rect 1782 -585 1787 -551
rect 1787 -585 1821 -551
rect 1821 -585 1834 -551
rect 1782 -592 1834 -585
rect 1846 -551 1898 -540
rect 1846 -585 1859 -551
rect 1859 -585 1893 -551
rect 1893 -585 1898 -551
rect 1846 -592 1898 -585
rect 1910 -551 1962 -540
rect 1974 -551 2026 -540
rect 2038 -551 2090 -540
rect 2102 -551 2154 -540
rect 2166 -551 2218 -540
rect 2230 -551 2282 -540
rect 2294 -551 2346 -540
rect 1910 -585 1931 -551
rect 1931 -585 1962 -551
rect 1974 -585 2003 -551
rect 2003 -585 2026 -551
rect 2038 -585 2075 -551
rect 2075 -585 2090 -551
rect 2102 -585 2109 -551
rect 2109 -585 2147 -551
rect 2147 -585 2154 -551
rect 2166 -585 2181 -551
rect 2181 -585 2218 -551
rect 2230 -585 2253 -551
rect 2253 -585 2282 -551
rect 2294 -585 2325 -551
rect 2325 -585 2346 -551
rect 1910 -592 1962 -585
rect 1974 -592 2026 -585
rect 2038 -592 2090 -585
rect 2102 -592 2154 -585
rect 2166 -592 2218 -585
rect 2230 -592 2282 -585
rect 2294 -592 2346 -585
rect 2358 -551 2410 -540
rect 2358 -585 2363 -551
rect 2363 -585 2397 -551
rect 2397 -585 2410 -551
rect 2358 -592 2410 -585
rect 2422 -551 2474 -540
rect 2422 -585 2435 -551
rect 2435 -585 2469 -551
rect 2469 -585 2474 -551
rect 2422 -592 2474 -585
rect 2486 -551 2538 -540
rect 2550 -551 2602 -540
rect 2614 -551 2666 -540
rect 2678 -551 2730 -540
rect 2742 -551 2794 -540
rect 2806 -551 2858 -540
rect 2870 -551 2922 -540
rect 2486 -585 2507 -551
rect 2507 -585 2538 -551
rect 2550 -585 2579 -551
rect 2579 -585 2602 -551
rect 2614 -585 2651 -551
rect 2651 -585 2666 -551
rect 2678 -585 2685 -551
rect 2685 -585 2723 -551
rect 2723 -585 2730 -551
rect 2742 -585 2757 -551
rect 2757 -585 2794 -551
rect 2806 -585 2829 -551
rect 2829 -585 2858 -551
rect 2870 -585 2901 -551
rect 2901 -585 2922 -551
rect 2486 -592 2538 -585
rect 2550 -592 2602 -585
rect 2614 -592 2666 -585
rect 2678 -592 2730 -585
rect 2742 -592 2794 -585
rect 2806 -592 2858 -585
rect 2870 -592 2922 -585
rect 2934 -551 2986 -540
rect 2934 -585 2939 -551
rect 2939 -585 2973 -551
rect 2973 -585 2986 -551
rect 2934 -592 2986 -585
rect 2998 -551 3050 -540
rect 2998 -585 3011 -551
rect 3011 -585 3045 -551
rect 3045 -585 3050 -551
rect 2998 -592 3050 -585
rect 3062 -551 3114 -540
rect 3126 -551 3178 -540
rect 3190 -551 3242 -540
rect 3254 -551 3306 -540
rect 3318 -551 3370 -540
rect 3382 -551 3434 -540
rect 3446 -551 3498 -540
rect 3062 -585 3083 -551
rect 3083 -585 3114 -551
rect 3126 -585 3155 -551
rect 3155 -585 3178 -551
rect 3190 -585 3227 -551
rect 3227 -585 3242 -551
rect 3254 -585 3261 -551
rect 3261 -585 3299 -551
rect 3299 -585 3306 -551
rect 3318 -585 3333 -551
rect 3333 -585 3370 -551
rect 3382 -585 3405 -551
rect 3405 -585 3434 -551
rect 3446 -585 3477 -551
rect 3477 -585 3498 -551
rect 3062 -592 3114 -585
rect 3126 -592 3178 -585
rect 3190 -592 3242 -585
rect 3254 -592 3306 -585
rect 3318 -592 3370 -585
rect 3382 -592 3434 -585
rect 3446 -592 3498 -585
rect 3510 -551 3562 -540
rect 3510 -585 3515 -551
rect 3515 -585 3549 -551
rect 3549 -585 3562 -551
rect 3510 -592 3562 -585
rect 3574 -551 3626 -540
rect 3574 -585 3587 -551
rect 3587 -585 3621 -551
rect 3621 -585 3626 -551
rect 3574 -592 3626 -585
rect 3638 -551 3690 -540
rect 3702 -551 3754 -540
rect 3766 -551 3818 -540
rect 3830 -551 3882 -540
rect 3894 -551 3946 -540
rect 3958 -551 4010 -540
rect 4022 -551 4074 -540
rect 3638 -585 3659 -551
rect 3659 -585 3690 -551
rect 3702 -585 3731 -551
rect 3731 -585 3754 -551
rect 3766 -585 3803 -551
rect 3803 -585 3818 -551
rect 3830 -585 3837 -551
rect 3837 -585 3875 -551
rect 3875 -585 3882 -551
rect 3894 -585 3909 -551
rect 3909 -585 3946 -551
rect 3958 -585 3981 -551
rect 3981 -585 4010 -551
rect 4022 -585 4053 -551
rect 4053 -585 4074 -551
rect 3638 -592 3690 -585
rect 3702 -592 3754 -585
rect 3766 -592 3818 -585
rect 3830 -592 3882 -585
rect 3894 -592 3946 -585
rect 3958 -592 4010 -585
rect 4022 -592 4074 -585
rect 4086 -551 4138 -540
rect 4086 -585 4091 -551
rect 4091 -585 4125 -551
rect 4125 -585 4138 -551
rect 4086 -592 4138 -585
rect 90 -817 142 -765
rect 90 -881 142 -829
rect 90 -945 142 -893
rect 90 -1009 142 -957
rect 282 -817 334 -765
rect 282 -881 334 -829
rect 282 -945 334 -893
rect 282 -1009 334 -957
rect 474 -817 526 -765
rect 474 -881 526 -829
rect 474 -945 526 -893
rect 474 -1009 526 -957
rect 666 -817 718 -765
rect 666 -881 718 -829
rect 666 -945 718 -893
rect 666 -1009 718 -957
rect 858 -817 910 -765
rect 858 -881 910 -829
rect 858 -945 910 -893
rect 858 -1009 910 -957
rect 1050 -817 1102 -765
rect 1050 -881 1102 -829
rect 1050 -945 1102 -893
rect 1050 -1009 1102 -957
rect 1242 -817 1294 -765
rect 1242 -881 1294 -829
rect 1242 -945 1294 -893
rect 1242 -1009 1294 -957
rect 1434 -817 1486 -765
rect 1434 -881 1486 -829
rect 1434 -945 1486 -893
rect 1434 -1009 1486 -957
rect 1626 -817 1678 -765
rect 1626 -881 1678 -829
rect 1626 -945 1678 -893
rect 1626 -1009 1678 -957
rect 1818 -817 1870 -765
rect 1818 -881 1870 -829
rect 1818 -945 1870 -893
rect 1818 -1009 1870 -957
rect 2010 -817 2062 -765
rect 2010 -881 2062 -829
rect 2010 -945 2062 -893
rect 2010 -1009 2062 -957
rect 2202 -817 2254 -765
rect 2202 -881 2254 -829
rect 2202 -945 2254 -893
rect 2202 -1009 2254 -957
rect 2394 -817 2446 -765
rect 2394 -881 2446 -829
rect 2394 -945 2446 -893
rect 2394 -1009 2446 -957
rect 2586 -817 2638 -765
rect 2586 -881 2638 -829
rect 2586 -945 2638 -893
rect 2586 -1009 2638 -957
rect 2778 -817 2830 -765
rect 2778 -881 2830 -829
rect 2778 -945 2830 -893
rect 2778 -1009 2830 -957
rect 2970 -817 3022 -765
rect 2970 -881 3022 -829
rect 2970 -945 3022 -893
rect 2970 -1009 3022 -957
rect 3162 -817 3214 -765
rect 3162 -881 3214 -829
rect 3162 -945 3214 -893
rect 3162 -1009 3214 -957
rect 3354 -817 3406 -765
rect 3354 -881 3406 -829
rect 3354 -945 3406 -893
rect 3354 -1009 3406 -957
rect 3546 -817 3598 -765
rect 3546 -881 3598 -829
rect 3546 -945 3598 -893
rect 3546 -1009 3598 -957
rect 3738 -817 3790 -765
rect 3738 -881 3790 -829
rect 3738 -945 3790 -893
rect 3738 -1009 3790 -957
rect 3930 -817 3982 -765
rect 3930 -881 3982 -829
rect 3930 -945 3982 -893
rect 3930 -1009 3982 -957
rect 4122 -817 4174 -765
rect 4122 -881 4174 -829
rect 4122 -945 4174 -893
rect 4122 -1009 4174 -957
rect 186 -1141 238 -1089
rect 186 -1205 238 -1153
rect 186 -1269 238 -1217
rect 186 -1333 238 -1281
rect 378 -1141 430 -1089
rect 378 -1205 430 -1153
rect 378 -1269 430 -1217
rect 378 -1333 430 -1281
rect 570 -1141 622 -1089
rect 570 -1205 622 -1153
rect 570 -1269 622 -1217
rect 570 -1333 622 -1281
rect 762 -1141 814 -1089
rect 762 -1205 814 -1153
rect 762 -1269 814 -1217
rect 762 -1333 814 -1281
rect 954 -1141 1006 -1089
rect 954 -1205 1006 -1153
rect 954 -1269 1006 -1217
rect 954 -1333 1006 -1281
rect 1146 -1141 1198 -1089
rect 1146 -1205 1198 -1153
rect 1146 -1269 1198 -1217
rect 1146 -1333 1198 -1281
rect 1338 -1141 1390 -1089
rect 1338 -1205 1390 -1153
rect 1338 -1269 1390 -1217
rect 1338 -1333 1390 -1281
rect 1530 -1141 1582 -1089
rect 1530 -1205 1582 -1153
rect 1530 -1269 1582 -1217
rect 1530 -1333 1582 -1281
rect 1722 -1141 1774 -1089
rect 1722 -1205 1774 -1153
rect 1722 -1269 1774 -1217
rect 1722 -1333 1774 -1281
rect 1914 -1141 1966 -1089
rect 1914 -1205 1966 -1153
rect 1914 -1269 1966 -1217
rect 1914 -1333 1966 -1281
rect 2106 -1141 2158 -1089
rect 2106 -1205 2158 -1153
rect 2106 -1269 2158 -1217
rect 2106 -1333 2158 -1281
rect 2298 -1141 2350 -1089
rect 2298 -1205 2350 -1153
rect 2298 -1269 2350 -1217
rect 2298 -1333 2350 -1281
rect 2490 -1141 2542 -1089
rect 2490 -1205 2542 -1153
rect 2490 -1269 2542 -1217
rect 2490 -1333 2542 -1281
rect 2682 -1141 2734 -1089
rect 2682 -1205 2734 -1153
rect 2682 -1269 2734 -1217
rect 2682 -1333 2734 -1281
rect 2874 -1141 2926 -1089
rect 2874 -1205 2926 -1153
rect 2874 -1269 2926 -1217
rect 2874 -1333 2926 -1281
rect 3066 -1141 3118 -1089
rect 3066 -1205 3118 -1153
rect 3066 -1269 3118 -1217
rect 3066 -1333 3118 -1281
rect 3258 -1141 3310 -1089
rect 3258 -1205 3310 -1153
rect 3258 -1269 3310 -1217
rect 3258 -1333 3310 -1281
rect 3450 -1141 3502 -1089
rect 3450 -1205 3502 -1153
rect 3450 -1269 3502 -1217
rect 3450 -1333 3502 -1281
rect 3642 -1141 3694 -1089
rect 3642 -1205 3694 -1153
rect 3642 -1269 3694 -1217
rect 3642 -1333 3694 -1281
rect 3834 -1141 3886 -1089
rect 3834 -1205 3886 -1153
rect 3834 -1269 3886 -1217
rect 3834 -1333 3886 -1281
rect 4026 -1141 4078 -1089
rect 4026 -1205 4078 -1153
rect 4026 -1269 4078 -1217
rect 4026 -1333 4078 -1281
<< metal2 >>
rect 82 -540 4182 -516
rect 82 -592 118 -540
rect 170 -592 182 -540
rect 234 -592 246 -540
rect 298 -592 310 -540
rect 362 -592 374 -540
rect 426 -592 438 -540
rect 490 -592 502 -540
rect 554 -592 566 -540
rect 618 -592 630 -540
rect 682 -592 694 -540
rect 746 -592 758 -540
rect 810 -592 822 -540
rect 874 -592 886 -540
rect 938 -592 950 -540
rect 1002 -592 1014 -540
rect 1066 -592 1078 -540
rect 1130 -592 1142 -540
rect 1194 -592 1206 -540
rect 1258 -592 1270 -540
rect 1322 -592 1334 -540
rect 1386 -592 1398 -540
rect 1450 -592 1462 -540
rect 1514 -592 1526 -540
rect 1578 -592 1590 -540
rect 1642 -592 1654 -540
rect 1706 -592 1718 -540
rect 1770 -592 1782 -540
rect 1834 -592 1846 -540
rect 1898 -592 1910 -540
rect 1962 -592 1974 -540
rect 2026 -592 2038 -540
rect 2090 -592 2102 -540
rect 2154 -592 2166 -540
rect 2218 -592 2230 -540
rect 2282 -592 2294 -540
rect 2346 -592 2358 -540
rect 2410 -592 2422 -540
rect 2474 -592 2486 -540
rect 2538 -592 2550 -540
rect 2602 -592 2614 -540
rect 2666 -592 2678 -540
rect 2730 -592 2742 -540
rect 2794 -592 2806 -540
rect 2858 -592 2870 -540
rect 2922 -592 2934 -540
rect 2986 -592 2998 -540
rect 3050 -592 3062 -540
rect 3114 -592 3126 -540
rect 3178 -592 3190 -540
rect 3242 -592 3254 -540
rect 3306 -592 3318 -540
rect 3370 -592 3382 -540
rect 3434 -592 3446 -540
rect 3498 -592 3510 -540
rect 3562 -592 3574 -540
rect 3626 -592 3638 -540
rect 3690 -592 3702 -540
rect 3754 -592 3766 -540
rect 3818 -592 3830 -540
rect 3882 -592 3894 -540
rect 3946 -592 3958 -540
rect 4010 -592 4022 -540
rect 4074 -592 4086 -540
rect 4138 -592 4182 -540
rect 82 -622 4182 -592
rect 82 -765 150 -622
rect 82 -817 90 -765
rect 142 -817 150 -765
rect 82 -829 150 -817
rect 82 -881 90 -829
rect 142 -881 150 -829
rect 82 -893 150 -881
rect 82 -945 90 -893
rect 142 -945 150 -893
rect 82 -957 150 -945
rect 82 -1009 90 -957
rect 142 -1009 150 -957
rect 82 -1032 150 -1009
rect 274 -765 342 -622
rect 274 -817 282 -765
rect 334 -817 342 -765
rect 274 -829 342 -817
rect 274 -881 282 -829
rect 334 -881 342 -829
rect 274 -893 342 -881
rect 274 -945 282 -893
rect 334 -945 342 -893
rect 274 -957 342 -945
rect 274 -1009 282 -957
rect 334 -1009 342 -957
rect 274 -1032 342 -1009
rect 466 -765 534 -622
rect 466 -817 474 -765
rect 526 -817 534 -765
rect 466 -829 534 -817
rect 466 -881 474 -829
rect 526 -881 534 -829
rect 466 -893 534 -881
rect 466 -945 474 -893
rect 526 -945 534 -893
rect 466 -957 534 -945
rect 466 -1009 474 -957
rect 526 -1009 534 -957
rect 466 -1032 534 -1009
rect 658 -765 726 -622
rect 658 -817 666 -765
rect 718 -817 726 -765
rect 658 -829 726 -817
rect 658 -881 666 -829
rect 718 -881 726 -829
rect 658 -893 726 -881
rect 658 -945 666 -893
rect 718 -945 726 -893
rect 658 -957 726 -945
rect 658 -1009 666 -957
rect 718 -1009 726 -957
rect 658 -1032 726 -1009
rect 850 -765 918 -622
rect 850 -817 858 -765
rect 910 -817 918 -765
rect 850 -829 918 -817
rect 850 -881 858 -829
rect 910 -881 918 -829
rect 850 -893 918 -881
rect 850 -945 858 -893
rect 910 -945 918 -893
rect 850 -957 918 -945
rect 850 -1009 858 -957
rect 910 -1009 918 -957
rect 850 -1032 918 -1009
rect 1042 -765 1110 -622
rect 1042 -817 1050 -765
rect 1102 -817 1110 -765
rect 1042 -829 1110 -817
rect 1042 -881 1050 -829
rect 1102 -881 1110 -829
rect 1042 -893 1110 -881
rect 1042 -945 1050 -893
rect 1102 -945 1110 -893
rect 1042 -957 1110 -945
rect 1042 -1009 1050 -957
rect 1102 -1009 1110 -957
rect 1042 -1032 1110 -1009
rect 1234 -765 1302 -622
rect 1234 -817 1242 -765
rect 1294 -817 1302 -765
rect 1234 -829 1302 -817
rect 1234 -881 1242 -829
rect 1294 -881 1302 -829
rect 1234 -893 1302 -881
rect 1234 -945 1242 -893
rect 1294 -945 1302 -893
rect 1234 -957 1302 -945
rect 1234 -1009 1242 -957
rect 1294 -1009 1302 -957
rect 1234 -1032 1302 -1009
rect 1426 -765 1494 -622
rect 1426 -817 1434 -765
rect 1486 -817 1494 -765
rect 1426 -829 1494 -817
rect 1426 -881 1434 -829
rect 1486 -881 1494 -829
rect 1426 -893 1494 -881
rect 1426 -945 1434 -893
rect 1486 -945 1494 -893
rect 1426 -957 1494 -945
rect 1426 -1009 1434 -957
rect 1486 -1009 1494 -957
rect 1426 -1032 1494 -1009
rect 1618 -765 1686 -622
rect 1618 -817 1626 -765
rect 1678 -817 1686 -765
rect 1618 -829 1686 -817
rect 1618 -881 1626 -829
rect 1678 -881 1686 -829
rect 1618 -893 1686 -881
rect 1618 -945 1626 -893
rect 1678 -945 1686 -893
rect 1618 -957 1686 -945
rect 1618 -1009 1626 -957
rect 1678 -1009 1686 -957
rect 1618 -1032 1686 -1009
rect 1810 -765 1878 -622
rect 1810 -817 1818 -765
rect 1870 -817 1878 -765
rect 1810 -829 1878 -817
rect 1810 -881 1818 -829
rect 1870 -881 1878 -829
rect 1810 -893 1878 -881
rect 1810 -945 1818 -893
rect 1870 -945 1878 -893
rect 1810 -957 1878 -945
rect 1810 -1009 1818 -957
rect 1870 -1009 1878 -957
rect 1810 -1032 1878 -1009
rect 2002 -765 2070 -622
rect 2002 -817 2010 -765
rect 2062 -817 2070 -765
rect 2002 -829 2070 -817
rect 2002 -881 2010 -829
rect 2062 -881 2070 -829
rect 2002 -893 2070 -881
rect 2002 -945 2010 -893
rect 2062 -945 2070 -893
rect 2002 -957 2070 -945
rect 2002 -1009 2010 -957
rect 2062 -1009 2070 -957
rect 2002 -1032 2070 -1009
rect 2194 -765 2262 -622
rect 2194 -817 2202 -765
rect 2254 -817 2262 -765
rect 2194 -829 2262 -817
rect 2194 -881 2202 -829
rect 2254 -881 2262 -829
rect 2194 -893 2262 -881
rect 2194 -945 2202 -893
rect 2254 -945 2262 -893
rect 2194 -957 2262 -945
rect 2194 -1009 2202 -957
rect 2254 -1009 2262 -957
rect 2194 -1032 2262 -1009
rect 2386 -765 2454 -622
rect 2386 -817 2394 -765
rect 2446 -817 2454 -765
rect 2386 -829 2454 -817
rect 2386 -881 2394 -829
rect 2446 -881 2454 -829
rect 2386 -893 2454 -881
rect 2386 -945 2394 -893
rect 2446 -945 2454 -893
rect 2386 -957 2454 -945
rect 2386 -1009 2394 -957
rect 2446 -1009 2454 -957
rect 2386 -1032 2454 -1009
rect 2578 -765 2646 -622
rect 2578 -817 2586 -765
rect 2638 -817 2646 -765
rect 2578 -829 2646 -817
rect 2578 -881 2586 -829
rect 2638 -881 2646 -829
rect 2578 -893 2646 -881
rect 2578 -945 2586 -893
rect 2638 -945 2646 -893
rect 2578 -957 2646 -945
rect 2578 -1009 2586 -957
rect 2638 -1009 2646 -957
rect 2578 -1032 2646 -1009
rect 2770 -765 2838 -622
rect 2770 -817 2778 -765
rect 2830 -817 2838 -765
rect 2770 -829 2838 -817
rect 2770 -881 2778 -829
rect 2830 -881 2838 -829
rect 2770 -893 2838 -881
rect 2770 -945 2778 -893
rect 2830 -945 2838 -893
rect 2770 -957 2838 -945
rect 2770 -1009 2778 -957
rect 2830 -1009 2838 -957
rect 2770 -1032 2838 -1009
rect 2962 -765 3030 -622
rect 2962 -817 2970 -765
rect 3022 -817 3030 -765
rect 2962 -829 3030 -817
rect 2962 -881 2970 -829
rect 3022 -881 3030 -829
rect 2962 -893 3030 -881
rect 2962 -945 2970 -893
rect 3022 -945 3030 -893
rect 2962 -957 3030 -945
rect 2962 -1009 2970 -957
rect 3022 -1009 3030 -957
rect 2962 -1032 3030 -1009
rect 3154 -765 3222 -622
rect 3154 -817 3162 -765
rect 3214 -817 3222 -765
rect 3154 -829 3222 -817
rect 3154 -881 3162 -829
rect 3214 -881 3222 -829
rect 3154 -893 3222 -881
rect 3154 -945 3162 -893
rect 3214 -945 3222 -893
rect 3154 -957 3222 -945
rect 3154 -1009 3162 -957
rect 3214 -1009 3222 -957
rect 3154 -1032 3222 -1009
rect 3346 -765 3414 -622
rect 3346 -817 3354 -765
rect 3406 -817 3414 -765
rect 3346 -829 3414 -817
rect 3346 -881 3354 -829
rect 3406 -881 3414 -829
rect 3346 -893 3414 -881
rect 3346 -945 3354 -893
rect 3406 -945 3414 -893
rect 3346 -957 3414 -945
rect 3346 -1009 3354 -957
rect 3406 -1009 3414 -957
rect 3346 -1032 3414 -1009
rect 3538 -765 3606 -622
rect 3538 -817 3546 -765
rect 3598 -817 3606 -765
rect 3538 -829 3606 -817
rect 3538 -881 3546 -829
rect 3598 -881 3606 -829
rect 3538 -893 3606 -881
rect 3538 -945 3546 -893
rect 3598 -945 3606 -893
rect 3538 -957 3606 -945
rect 3538 -1009 3546 -957
rect 3598 -1009 3606 -957
rect 3538 -1032 3606 -1009
rect 3730 -765 3798 -622
rect 3730 -817 3738 -765
rect 3790 -817 3798 -765
rect 3730 -829 3798 -817
rect 3730 -881 3738 -829
rect 3790 -881 3798 -829
rect 3730 -893 3798 -881
rect 3730 -945 3738 -893
rect 3790 -945 3798 -893
rect 3730 -957 3798 -945
rect 3730 -1009 3738 -957
rect 3790 -1009 3798 -957
rect 3730 -1032 3798 -1009
rect 3922 -765 3990 -622
rect 3922 -817 3930 -765
rect 3982 -817 3990 -765
rect 3922 -829 3990 -817
rect 3922 -881 3930 -829
rect 3982 -881 3990 -829
rect 3922 -893 3990 -881
rect 3922 -945 3930 -893
rect 3982 -945 3990 -893
rect 3922 -957 3990 -945
rect 3922 -1009 3930 -957
rect 3982 -1009 3990 -957
rect 3922 -1032 3990 -1009
rect 4114 -765 4182 -622
rect 4114 -817 4122 -765
rect 4174 -817 4182 -765
rect 4114 -829 4182 -817
rect 4114 -881 4122 -829
rect 4174 -881 4182 -829
rect 4114 -893 4182 -881
rect 4114 -945 4122 -893
rect 4174 -945 4182 -893
rect 4114 -957 4182 -945
rect 4114 -1009 4122 -957
rect 4174 -1009 4182 -957
rect 4114 -1032 4182 -1009
rect 180 -1089 244 -1070
rect 180 -1102 186 -1089
rect 238 -1102 244 -1089
rect 180 -1158 184 -1102
rect 240 -1158 244 -1102
rect 180 -1182 186 -1158
rect 238 -1182 244 -1158
rect 180 -1238 184 -1182
rect 240 -1238 244 -1182
rect 180 -1262 186 -1238
rect 238 -1262 244 -1238
rect 180 -1318 184 -1262
rect 240 -1318 244 -1262
rect 180 -1333 186 -1318
rect 238 -1333 244 -1318
rect 180 -1350 244 -1333
rect 372 -1089 436 -1070
rect 372 -1102 378 -1089
rect 430 -1102 436 -1089
rect 372 -1158 376 -1102
rect 432 -1158 436 -1102
rect 372 -1182 378 -1158
rect 430 -1182 436 -1158
rect 372 -1238 376 -1182
rect 432 -1238 436 -1182
rect 372 -1262 378 -1238
rect 430 -1262 436 -1238
rect 372 -1318 376 -1262
rect 432 -1318 436 -1262
rect 372 -1333 378 -1318
rect 430 -1333 436 -1318
rect 372 -1350 436 -1333
rect 564 -1089 628 -1070
rect 564 -1102 570 -1089
rect 622 -1102 628 -1089
rect 564 -1158 568 -1102
rect 624 -1158 628 -1102
rect 564 -1182 570 -1158
rect 622 -1182 628 -1158
rect 564 -1238 568 -1182
rect 624 -1238 628 -1182
rect 564 -1262 570 -1238
rect 622 -1262 628 -1238
rect 564 -1318 568 -1262
rect 624 -1318 628 -1262
rect 564 -1333 570 -1318
rect 622 -1333 628 -1318
rect 564 -1350 628 -1333
rect 756 -1089 820 -1070
rect 756 -1102 762 -1089
rect 814 -1102 820 -1089
rect 756 -1158 760 -1102
rect 816 -1158 820 -1102
rect 756 -1182 762 -1158
rect 814 -1182 820 -1158
rect 756 -1238 760 -1182
rect 816 -1238 820 -1182
rect 756 -1262 762 -1238
rect 814 -1262 820 -1238
rect 756 -1318 760 -1262
rect 816 -1318 820 -1262
rect 756 -1333 762 -1318
rect 814 -1333 820 -1318
rect 756 -1350 820 -1333
rect 948 -1089 1012 -1070
rect 948 -1102 954 -1089
rect 1006 -1102 1012 -1089
rect 948 -1158 952 -1102
rect 1008 -1158 1012 -1102
rect 948 -1182 954 -1158
rect 1006 -1182 1012 -1158
rect 948 -1238 952 -1182
rect 1008 -1238 1012 -1182
rect 948 -1262 954 -1238
rect 1006 -1262 1012 -1238
rect 948 -1318 952 -1262
rect 1008 -1318 1012 -1262
rect 948 -1333 954 -1318
rect 1006 -1333 1012 -1318
rect 948 -1350 1012 -1333
rect 1140 -1089 1204 -1070
rect 1140 -1102 1146 -1089
rect 1198 -1102 1204 -1089
rect 1140 -1158 1144 -1102
rect 1200 -1158 1204 -1102
rect 1140 -1182 1146 -1158
rect 1198 -1182 1204 -1158
rect 1140 -1238 1144 -1182
rect 1200 -1238 1204 -1182
rect 1140 -1262 1146 -1238
rect 1198 -1262 1204 -1238
rect 1140 -1318 1144 -1262
rect 1200 -1318 1204 -1262
rect 1140 -1333 1146 -1318
rect 1198 -1333 1204 -1318
rect 1140 -1350 1204 -1333
rect 1332 -1089 1396 -1070
rect 1332 -1102 1338 -1089
rect 1390 -1102 1396 -1089
rect 1332 -1158 1336 -1102
rect 1392 -1158 1396 -1102
rect 1332 -1182 1338 -1158
rect 1390 -1182 1396 -1158
rect 1332 -1238 1336 -1182
rect 1392 -1238 1396 -1182
rect 1332 -1262 1338 -1238
rect 1390 -1262 1396 -1238
rect 1332 -1318 1336 -1262
rect 1392 -1318 1396 -1262
rect 1332 -1333 1338 -1318
rect 1390 -1333 1396 -1318
rect 1332 -1350 1396 -1333
rect 1524 -1089 1588 -1070
rect 1524 -1102 1530 -1089
rect 1582 -1102 1588 -1089
rect 1524 -1158 1528 -1102
rect 1584 -1158 1588 -1102
rect 1524 -1182 1530 -1158
rect 1582 -1182 1588 -1158
rect 1524 -1238 1528 -1182
rect 1584 -1238 1588 -1182
rect 1524 -1262 1530 -1238
rect 1582 -1262 1588 -1238
rect 1524 -1318 1528 -1262
rect 1584 -1318 1588 -1262
rect 1524 -1333 1530 -1318
rect 1582 -1333 1588 -1318
rect 1524 -1350 1588 -1333
rect 1716 -1089 1780 -1070
rect 1716 -1102 1722 -1089
rect 1774 -1102 1780 -1089
rect 1716 -1158 1720 -1102
rect 1776 -1158 1780 -1102
rect 1716 -1182 1722 -1158
rect 1774 -1182 1780 -1158
rect 1716 -1238 1720 -1182
rect 1776 -1238 1780 -1182
rect 1716 -1262 1722 -1238
rect 1774 -1262 1780 -1238
rect 1716 -1318 1720 -1262
rect 1776 -1318 1780 -1262
rect 1716 -1333 1722 -1318
rect 1774 -1333 1780 -1318
rect 1716 -1350 1780 -1333
rect 1908 -1089 1972 -1070
rect 1908 -1102 1914 -1089
rect 1966 -1102 1972 -1089
rect 1908 -1158 1912 -1102
rect 1968 -1158 1972 -1102
rect 1908 -1182 1914 -1158
rect 1966 -1182 1972 -1158
rect 1908 -1238 1912 -1182
rect 1968 -1238 1972 -1182
rect 1908 -1262 1914 -1238
rect 1966 -1262 1972 -1238
rect 1908 -1318 1912 -1262
rect 1968 -1318 1972 -1262
rect 1908 -1333 1914 -1318
rect 1966 -1333 1972 -1318
rect 1908 -1350 1972 -1333
rect 2100 -1089 2164 -1070
rect 2100 -1102 2106 -1089
rect 2158 -1102 2164 -1089
rect 2100 -1158 2104 -1102
rect 2160 -1158 2164 -1102
rect 2100 -1182 2106 -1158
rect 2158 -1182 2164 -1158
rect 2100 -1238 2104 -1182
rect 2160 -1238 2164 -1182
rect 2100 -1262 2106 -1238
rect 2158 -1262 2164 -1238
rect 2100 -1318 2104 -1262
rect 2160 -1318 2164 -1262
rect 2100 -1333 2106 -1318
rect 2158 -1333 2164 -1318
rect 2100 -1350 2164 -1333
rect 2292 -1089 2356 -1070
rect 2292 -1102 2298 -1089
rect 2350 -1102 2356 -1089
rect 2292 -1158 2296 -1102
rect 2352 -1158 2356 -1102
rect 2292 -1182 2298 -1158
rect 2350 -1182 2356 -1158
rect 2292 -1238 2296 -1182
rect 2352 -1238 2356 -1182
rect 2292 -1262 2298 -1238
rect 2350 -1262 2356 -1238
rect 2292 -1318 2296 -1262
rect 2352 -1318 2356 -1262
rect 2292 -1333 2298 -1318
rect 2350 -1333 2356 -1318
rect 2292 -1350 2356 -1333
rect 2484 -1089 2548 -1070
rect 2484 -1102 2490 -1089
rect 2542 -1102 2548 -1089
rect 2484 -1158 2488 -1102
rect 2544 -1158 2548 -1102
rect 2484 -1182 2490 -1158
rect 2542 -1182 2548 -1158
rect 2484 -1238 2488 -1182
rect 2544 -1238 2548 -1182
rect 2484 -1262 2490 -1238
rect 2542 -1262 2548 -1238
rect 2484 -1318 2488 -1262
rect 2544 -1318 2548 -1262
rect 2484 -1333 2490 -1318
rect 2542 -1333 2548 -1318
rect 2484 -1350 2548 -1333
rect 2676 -1089 2740 -1070
rect 2676 -1102 2682 -1089
rect 2734 -1102 2740 -1089
rect 2676 -1158 2680 -1102
rect 2736 -1158 2740 -1102
rect 2676 -1182 2682 -1158
rect 2734 -1182 2740 -1158
rect 2676 -1238 2680 -1182
rect 2736 -1238 2740 -1182
rect 2676 -1262 2682 -1238
rect 2734 -1262 2740 -1238
rect 2676 -1318 2680 -1262
rect 2736 -1318 2740 -1262
rect 2676 -1333 2682 -1318
rect 2734 -1333 2740 -1318
rect 2676 -1350 2740 -1333
rect 2868 -1089 2932 -1070
rect 2868 -1102 2874 -1089
rect 2926 -1102 2932 -1089
rect 2868 -1158 2872 -1102
rect 2928 -1158 2932 -1102
rect 2868 -1182 2874 -1158
rect 2926 -1182 2932 -1158
rect 2868 -1238 2872 -1182
rect 2928 -1238 2932 -1182
rect 2868 -1262 2874 -1238
rect 2926 -1262 2932 -1238
rect 2868 -1318 2872 -1262
rect 2928 -1318 2932 -1262
rect 2868 -1333 2874 -1318
rect 2926 -1333 2932 -1318
rect 2868 -1350 2932 -1333
rect 3060 -1089 3124 -1070
rect 3060 -1102 3066 -1089
rect 3118 -1102 3124 -1089
rect 3060 -1158 3064 -1102
rect 3120 -1158 3124 -1102
rect 3060 -1182 3066 -1158
rect 3118 -1182 3124 -1158
rect 3060 -1238 3064 -1182
rect 3120 -1238 3124 -1182
rect 3060 -1262 3066 -1238
rect 3118 -1262 3124 -1238
rect 3060 -1318 3064 -1262
rect 3120 -1318 3124 -1262
rect 3060 -1333 3066 -1318
rect 3118 -1333 3124 -1318
rect 3060 -1350 3124 -1333
rect 3252 -1089 3316 -1070
rect 3252 -1102 3258 -1089
rect 3310 -1102 3316 -1089
rect 3252 -1158 3256 -1102
rect 3312 -1158 3316 -1102
rect 3252 -1182 3258 -1158
rect 3310 -1182 3316 -1158
rect 3252 -1238 3256 -1182
rect 3312 -1238 3316 -1182
rect 3252 -1262 3258 -1238
rect 3310 -1262 3316 -1238
rect 3252 -1318 3256 -1262
rect 3312 -1318 3316 -1262
rect 3252 -1333 3258 -1318
rect 3310 -1333 3316 -1318
rect 3252 -1350 3316 -1333
rect 3444 -1089 3508 -1070
rect 3444 -1102 3450 -1089
rect 3502 -1102 3508 -1089
rect 3444 -1158 3448 -1102
rect 3504 -1158 3508 -1102
rect 3444 -1182 3450 -1158
rect 3502 -1182 3508 -1158
rect 3444 -1238 3448 -1182
rect 3504 -1238 3508 -1182
rect 3444 -1262 3450 -1238
rect 3502 -1262 3508 -1238
rect 3444 -1318 3448 -1262
rect 3504 -1318 3508 -1262
rect 3444 -1333 3450 -1318
rect 3502 -1333 3508 -1318
rect 3444 -1350 3508 -1333
rect 3636 -1089 3700 -1070
rect 3636 -1102 3642 -1089
rect 3694 -1102 3700 -1089
rect 3636 -1158 3640 -1102
rect 3696 -1158 3700 -1102
rect 3636 -1182 3642 -1158
rect 3694 -1182 3700 -1158
rect 3636 -1238 3640 -1182
rect 3696 -1238 3700 -1182
rect 3636 -1262 3642 -1238
rect 3694 -1262 3700 -1238
rect 3636 -1318 3640 -1262
rect 3696 -1318 3700 -1262
rect 3636 -1333 3642 -1318
rect 3694 -1333 3700 -1318
rect 3636 -1350 3700 -1333
rect 3828 -1089 3892 -1070
rect 3828 -1102 3834 -1089
rect 3886 -1102 3892 -1089
rect 3828 -1158 3832 -1102
rect 3888 -1158 3892 -1102
rect 3828 -1182 3834 -1158
rect 3886 -1182 3892 -1158
rect 3828 -1238 3832 -1182
rect 3888 -1238 3892 -1182
rect 3828 -1262 3834 -1238
rect 3886 -1262 3892 -1238
rect 3828 -1318 3832 -1262
rect 3888 -1318 3892 -1262
rect 3828 -1333 3834 -1318
rect 3886 -1333 3892 -1318
rect 3828 -1350 3892 -1333
rect 4020 -1089 4084 -1070
rect 4020 -1102 4026 -1089
rect 4078 -1102 4084 -1089
rect 4020 -1158 4024 -1102
rect 4080 -1158 4084 -1102
rect 4020 -1182 4026 -1158
rect 4078 -1182 4084 -1158
rect 4020 -1238 4024 -1182
rect 4080 -1238 4084 -1182
rect 4020 -1262 4026 -1238
rect 4078 -1262 4084 -1238
rect 4020 -1318 4024 -1262
rect 4080 -1318 4084 -1262
rect 4020 -1333 4026 -1318
rect 4078 -1333 4084 -1318
rect 4020 -1350 4084 -1333
<< via2 >>
rect 184 -1141 186 -1102
rect 186 -1141 238 -1102
rect 238 -1141 240 -1102
rect 184 -1153 240 -1141
rect 184 -1158 186 -1153
rect 186 -1158 238 -1153
rect 238 -1158 240 -1153
rect 184 -1205 186 -1182
rect 186 -1205 238 -1182
rect 238 -1205 240 -1182
rect 184 -1217 240 -1205
rect 184 -1238 186 -1217
rect 186 -1238 238 -1217
rect 238 -1238 240 -1217
rect 184 -1269 186 -1262
rect 186 -1269 238 -1262
rect 238 -1269 240 -1262
rect 184 -1281 240 -1269
rect 184 -1318 186 -1281
rect 186 -1318 238 -1281
rect 238 -1318 240 -1281
rect 376 -1141 378 -1102
rect 378 -1141 430 -1102
rect 430 -1141 432 -1102
rect 376 -1153 432 -1141
rect 376 -1158 378 -1153
rect 378 -1158 430 -1153
rect 430 -1158 432 -1153
rect 376 -1205 378 -1182
rect 378 -1205 430 -1182
rect 430 -1205 432 -1182
rect 376 -1217 432 -1205
rect 376 -1238 378 -1217
rect 378 -1238 430 -1217
rect 430 -1238 432 -1217
rect 376 -1269 378 -1262
rect 378 -1269 430 -1262
rect 430 -1269 432 -1262
rect 376 -1281 432 -1269
rect 376 -1318 378 -1281
rect 378 -1318 430 -1281
rect 430 -1318 432 -1281
rect 568 -1141 570 -1102
rect 570 -1141 622 -1102
rect 622 -1141 624 -1102
rect 568 -1153 624 -1141
rect 568 -1158 570 -1153
rect 570 -1158 622 -1153
rect 622 -1158 624 -1153
rect 568 -1205 570 -1182
rect 570 -1205 622 -1182
rect 622 -1205 624 -1182
rect 568 -1217 624 -1205
rect 568 -1238 570 -1217
rect 570 -1238 622 -1217
rect 622 -1238 624 -1217
rect 568 -1269 570 -1262
rect 570 -1269 622 -1262
rect 622 -1269 624 -1262
rect 568 -1281 624 -1269
rect 568 -1318 570 -1281
rect 570 -1318 622 -1281
rect 622 -1318 624 -1281
rect 760 -1141 762 -1102
rect 762 -1141 814 -1102
rect 814 -1141 816 -1102
rect 760 -1153 816 -1141
rect 760 -1158 762 -1153
rect 762 -1158 814 -1153
rect 814 -1158 816 -1153
rect 760 -1205 762 -1182
rect 762 -1205 814 -1182
rect 814 -1205 816 -1182
rect 760 -1217 816 -1205
rect 760 -1238 762 -1217
rect 762 -1238 814 -1217
rect 814 -1238 816 -1217
rect 760 -1269 762 -1262
rect 762 -1269 814 -1262
rect 814 -1269 816 -1262
rect 760 -1281 816 -1269
rect 760 -1318 762 -1281
rect 762 -1318 814 -1281
rect 814 -1318 816 -1281
rect 952 -1141 954 -1102
rect 954 -1141 1006 -1102
rect 1006 -1141 1008 -1102
rect 952 -1153 1008 -1141
rect 952 -1158 954 -1153
rect 954 -1158 1006 -1153
rect 1006 -1158 1008 -1153
rect 952 -1205 954 -1182
rect 954 -1205 1006 -1182
rect 1006 -1205 1008 -1182
rect 952 -1217 1008 -1205
rect 952 -1238 954 -1217
rect 954 -1238 1006 -1217
rect 1006 -1238 1008 -1217
rect 952 -1269 954 -1262
rect 954 -1269 1006 -1262
rect 1006 -1269 1008 -1262
rect 952 -1281 1008 -1269
rect 952 -1318 954 -1281
rect 954 -1318 1006 -1281
rect 1006 -1318 1008 -1281
rect 1144 -1141 1146 -1102
rect 1146 -1141 1198 -1102
rect 1198 -1141 1200 -1102
rect 1144 -1153 1200 -1141
rect 1144 -1158 1146 -1153
rect 1146 -1158 1198 -1153
rect 1198 -1158 1200 -1153
rect 1144 -1205 1146 -1182
rect 1146 -1205 1198 -1182
rect 1198 -1205 1200 -1182
rect 1144 -1217 1200 -1205
rect 1144 -1238 1146 -1217
rect 1146 -1238 1198 -1217
rect 1198 -1238 1200 -1217
rect 1144 -1269 1146 -1262
rect 1146 -1269 1198 -1262
rect 1198 -1269 1200 -1262
rect 1144 -1281 1200 -1269
rect 1144 -1318 1146 -1281
rect 1146 -1318 1198 -1281
rect 1198 -1318 1200 -1281
rect 1336 -1141 1338 -1102
rect 1338 -1141 1390 -1102
rect 1390 -1141 1392 -1102
rect 1336 -1153 1392 -1141
rect 1336 -1158 1338 -1153
rect 1338 -1158 1390 -1153
rect 1390 -1158 1392 -1153
rect 1336 -1205 1338 -1182
rect 1338 -1205 1390 -1182
rect 1390 -1205 1392 -1182
rect 1336 -1217 1392 -1205
rect 1336 -1238 1338 -1217
rect 1338 -1238 1390 -1217
rect 1390 -1238 1392 -1217
rect 1336 -1269 1338 -1262
rect 1338 -1269 1390 -1262
rect 1390 -1269 1392 -1262
rect 1336 -1281 1392 -1269
rect 1336 -1318 1338 -1281
rect 1338 -1318 1390 -1281
rect 1390 -1318 1392 -1281
rect 1528 -1141 1530 -1102
rect 1530 -1141 1582 -1102
rect 1582 -1141 1584 -1102
rect 1528 -1153 1584 -1141
rect 1528 -1158 1530 -1153
rect 1530 -1158 1582 -1153
rect 1582 -1158 1584 -1153
rect 1528 -1205 1530 -1182
rect 1530 -1205 1582 -1182
rect 1582 -1205 1584 -1182
rect 1528 -1217 1584 -1205
rect 1528 -1238 1530 -1217
rect 1530 -1238 1582 -1217
rect 1582 -1238 1584 -1217
rect 1528 -1269 1530 -1262
rect 1530 -1269 1582 -1262
rect 1582 -1269 1584 -1262
rect 1528 -1281 1584 -1269
rect 1528 -1318 1530 -1281
rect 1530 -1318 1582 -1281
rect 1582 -1318 1584 -1281
rect 1720 -1141 1722 -1102
rect 1722 -1141 1774 -1102
rect 1774 -1141 1776 -1102
rect 1720 -1153 1776 -1141
rect 1720 -1158 1722 -1153
rect 1722 -1158 1774 -1153
rect 1774 -1158 1776 -1153
rect 1720 -1205 1722 -1182
rect 1722 -1205 1774 -1182
rect 1774 -1205 1776 -1182
rect 1720 -1217 1776 -1205
rect 1720 -1238 1722 -1217
rect 1722 -1238 1774 -1217
rect 1774 -1238 1776 -1217
rect 1720 -1269 1722 -1262
rect 1722 -1269 1774 -1262
rect 1774 -1269 1776 -1262
rect 1720 -1281 1776 -1269
rect 1720 -1318 1722 -1281
rect 1722 -1318 1774 -1281
rect 1774 -1318 1776 -1281
rect 1912 -1141 1914 -1102
rect 1914 -1141 1966 -1102
rect 1966 -1141 1968 -1102
rect 1912 -1153 1968 -1141
rect 1912 -1158 1914 -1153
rect 1914 -1158 1966 -1153
rect 1966 -1158 1968 -1153
rect 1912 -1205 1914 -1182
rect 1914 -1205 1966 -1182
rect 1966 -1205 1968 -1182
rect 1912 -1217 1968 -1205
rect 1912 -1238 1914 -1217
rect 1914 -1238 1966 -1217
rect 1966 -1238 1968 -1217
rect 1912 -1269 1914 -1262
rect 1914 -1269 1966 -1262
rect 1966 -1269 1968 -1262
rect 1912 -1281 1968 -1269
rect 1912 -1318 1914 -1281
rect 1914 -1318 1966 -1281
rect 1966 -1318 1968 -1281
rect 2104 -1141 2106 -1102
rect 2106 -1141 2158 -1102
rect 2158 -1141 2160 -1102
rect 2104 -1153 2160 -1141
rect 2104 -1158 2106 -1153
rect 2106 -1158 2158 -1153
rect 2158 -1158 2160 -1153
rect 2104 -1205 2106 -1182
rect 2106 -1205 2158 -1182
rect 2158 -1205 2160 -1182
rect 2104 -1217 2160 -1205
rect 2104 -1238 2106 -1217
rect 2106 -1238 2158 -1217
rect 2158 -1238 2160 -1217
rect 2104 -1269 2106 -1262
rect 2106 -1269 2158 -1262
rect 2158 -1269 2160 -1262
rect 2104 -1281 2160 -1269
rect 2104 -1318 2106 -1281
rect 2106 -1318 2158 -1281
rect 2158 -1318 2160 -1281
rect 2296 -1141 2298 -1102
rect 2298 -1141 2350 -1102
rect 2350 -1141 2352 -1102
rect 2296 -1153 2352 -1141
rect 2296 -1158 2298 -1153
rect 2298 -1158 2350 -1153
rect 2350 -1158 2352 -1153
rect 2296 -1205 2298 -1182
rect 2298 -1205 2350 -1182
rect 2350 -1205 2352 -1182
rect 2296 -1217 2352 -1205
rect 2296 -1238 2298 -1217
rect 2298 -1238 2350 -1217
rect 2350 -1238 2352 -1217
rect 2296 -1269 2298 -1262
rect 2298 -1269 2350 -1262
rect 2350 -1269 2352 -1262
rect 2296 -1281 2352 -1269
rect 2296 -1318 2298 -1281
rect 2298 -1318 2350 -1281
rect 2350 -1318 2352 -1281
rect 2488 -1141 2490 -1102
rect 2490 -1141 2542 -1102
rect 2542 -1141 2544 -1102
rect 2488 -1153 2544 -1141
rect 2488 -1158 2490 -1153
rect 2490 -1158 2542 -1153
rect 2542 -1158 2544 -1153
rect 2488 -1205 2490 -1182
rect 2490 -1205 2542 -1182
rect 2542 -1205 2544 -1182
rect 2488 -1217 2544 -1205
rect 2488 -1238 2490 -1217
rect 2490 -1238 2542 -1217
rect 2542 -1238 2544 -1217
rect 2488 -1269 2490 -1262
rect 2490 -1269 2542 -1262
rect 2542 -1269 2544 -1262
rect 2488 -1281 2544 -1269
rect 2488 -1318 2490 -1281
rect 2490 -1318 2542 -1281
rect 2542 -1318 2544 -1281
rect 2680 -1141 2682 -1102
rect 2682 -1141 2734 -1102
rect 2734 -1141 2736 -1102
rect 2680 -1153 2736 -1141
rect 2680 -1158 2682 -1153
rect 2682 -1158 2734 -1153
rect 2734 -1158 2736 -1153
rect 2680 -1205 2682 -1182
rect 2682 -1205 2734 -1182
rect 2734 -1205 2736 -1182
rect 2680 -1217 2736 -1205
rect 2680 -1238 2682 -1217
rect 2682 -1238 2734 -1217
rect 2734 -1238 2736 -1217
rect 2680 -1269 2682 -1262
rect 2682 -1269 2734 -1262
rect 2734 -1269 2736 -1262
rect 2680 -1281 2736 -1269
rect 2680 -1318 2682 -1281
rect 2682 -1318 2734 -1281
rect 2734 -1318 2736 -1281
rect 2872 -1141 2874 -1102
rect 2874 -1141 2926 -1102
rect 2926 -1141 2928 -1102
rect 2872 -1153 2928 -1141
rect 2872 -1158 2874 -1153
rect 2874 -1158 2926 -1153
rect 2926 -1158 2928 -1153
rect 2872 -1205 2874 -1182
rect 2874 -1205 2926 -1182
rect 2926 -1205 2928 -1182
rect 2872 -1217 2928 -1205
rect 2872 -1238 2874 -1217
rect 2874 -1238 2926 -1217
rect 2926 -1238 2928 -1217
rect 2872 -1269 2874 -1262
rect 2874 -1269 2926 -1262
rect 2926 -1269 2928 -1262
rect 2872 -1281 2928 -1269
rect 2872 -1318 2874 -1281
rect 2874 -1318 2926 -1281
rect 2926 -1318 2928 -1281
rect 3064 -1141 3066 -1102
rect 3066 -1141 3118 -1102
rect 3118 -1141 3120 -1102
rect 3064 -1153 3120 -1141
rect 3064 -1158 3066 -1153
rect 3066 -1158 3118 -1153
rect 3118 -1158 3120 -1153
rect 3064 -1205 3066 -1182
rect 3066 -1205 3118 -1182
rect 3118 -1205 3120 -1182
rect 3064 -1217 3120 -1205
rect 3064 -1238 3066 -1217
rect 3066 -1238 3118 -1217
rect 3118 -1238 3120 -1217
rect 3064 -1269 3066 -1262
rect 3066 -1269 3118 -1262
rect 3118 -1269 3120 -1262
rect 3064 -1281 3120 -1269
rect 3064 -1318 3066 -1281
rect 3066 -1318 3118 -1281
rect 3118 -1318 3120 -1281
rect 3256 -1141 3258 -1102
rect 3258 -1141 3310 -1102
rect 3310 -1141 3312 -1102
rect 3256 -1153 3312 -1141
rect 3256 -1158 3258 -1153
rect 3258 -1158 3310 -1153
rect 3310 -1158 3312 -1153
rect 3256 -1205 3258 -1182
rect 3258 -1205 3310 -1182
rect 3310 -1205 3312 -1182
rect 3256 -1217 3312 -1205
rect 3256 -1238 3258 -1217
rect 3258 -1238 3310 -1217
rect 3310 -1238 3312 -1217
rect 3256 -1269 3258 -1262
rect 3258 -1269 3310 -1262
rect 3310 -1269 3312 -1262
rect 3256 -1281 3312 -1269
rect 3256 -1318 3258 -1281
rect 3258 -1318 3310 -1281
rect 3310 -1318 3312 -1281
rect 3448 -1141 3450 -1102
rect 3450 -1141 3502 -1102
rect 3502 -1141 3504 -1102
rect 3448 -1153 3504 -1141
rect 3448 -1158 3450 -1153
rect 3450 -1158 3502 -1153
rect 3502 -1158 3504 -1153
rect 3448 -1205 3450 -1182
rect 3450 -1205 3502 -1182
rect 3502 -1205 3504 -1182
rect 3448 -1217 3504 -1205
rect 3448 -1238 3450 -1217
rect 3450 -1238 3502 -1217
rect 3502 -1238 3504 -1217
rect 3448 -1269 3450 -1262
rect 3450 -1269 3502 -1262
rect 3502 -1269 3504 -1262
rect 3448 -1281 3504 -1269
rect 3448 -1318 3450 -1281
rect 3450 -1318 3502 -1281
rect 3502 -1318 3504 -1281
rect 3640 -1141 3642 -1102
rect 3642 -1141 3694 -1102
rect 3694 -1141 3696 -1102
rect 3640 -1153 3696 -1141
rect 3640 -1158 3642 -1153
rect 3642 -1158 3694 -1153
rect 3694 -1158 3696 -1153
rect 3640 -1205 3642 -1182
rect 3642 -1205 3694 -1182
rect 3694 -1205 3696 -1182
rect 3640 -1217 3696 -1205
rect 3640 -1238 3642 -1217
rect 3642 -1238 3694 -1217
rect 3694 -1238 3696 -1217
rect 3640 -1269 3642 -1262
rect 3642 -1269 3694 -1262
rect 3694 -1269 3696 -1262
rect 3640 -1281 3696 -1269
rect 3640 -1318 3642 -1281
rect 3642 -1318 3694 -1281
rect 3694 -1318 3696 -1281
rect 3832 -1141 3834 -1102
rect 3834 -1141 3886 -1102
rect 3886 -1141 3888 -1102
rect 3832 -1153 3888 -1141
rect 3832 -1158 3834 -1153
rect 3834 -1158 3886 -1153
rect 3886 -1158 3888 -1153
rect 3832 -1205 3834 -1182
rect 3834 -1205 3886 -1182
rect 3886 -1205 3888 -1182
rect 3832 -1217 3888 -1205
rect 3832 -1238 3834 -1217
rect 3834 -1238 3886 -1217
rect 3886 -1238 3888 -1217
rect 3832 -1269 3834 -1262
rect 3834 -1269 3886 -1262
rect 3886 -1269 3888 -1262
rect 3832 -1281 3888 -1269
rect 3832 -1318 3834 -1281
rect 3834 -1318 3886 -1281
rect 3886 -1318 3888 -1281
rect 4024 -1141 4026 -1102
rect 4026 -1141 4078 -1102
rect 4078 -1141 4080 -1102
rect 4024 -1153 4080 -1141
rect 4024 -1158 4026 -1153
rect 4026 -1158 4078 -1153
rect 4078 -1158 4080 -1153
rect 4024 -1205 4026 -1182
rect 4026 -1205 4078 -1182
rect 4078 -1205 4080 -1182
rect 4024 -1217 4080 -1205
rect 4024 -1238 4026 -1217
rect 4026 -1238 4078 -1217
rect 4078 -1238 4080 -1217
rect 4024 -1269 4026 -1262
rect 4026 -1269 4078 -1262
rect 4078 -1269 4080 -1262
rect 4024 -1281 4080 -1269
rect 4024 -1318 4026 -1281
rect 4026 -1318 4078 -1281
rect 4078 -1318 4080 -1281
<< metal3 >>
rect 178 -1102 246 -1070
rect 178 -1158 184 -1102
rect 240 -1158 246 -1102
rect 178 -1182 246 -1158
rect 178 -1238 184 -1182
rect 240 -1238 246 -1182
rect 178 -1262 246 -1238
rect 178 -1318 184 -1262
rect 240 -1318 246 -1262
rect 178 -1396 246 -1318
rect 370 -1102 438 -1070
rect 370 -1158 376 -1102
rect 432 -1158 438 -1102
rect 370 -1182 438 -1158
rect 370 -1238 376 -1182
rect 432 -1238 438 -1182
rect 370 -1262 438 -1238
rect 370 -1318 376 -1262
rect 432 -1318 438 -1262
rect 370 -1396 438 -1318
rect 562 -1102 630 -1070
rect 562 -1158 568 -1102
rect 624 -1158 630 -1102
rect 562 -1182 630 -1158
rect 562 -1238 568 -1182
rect 624 -1238 630 -1182
rect 562 -1262 630 -1238
rect 562 -1318 568 -1262
rect 624 -1318 630 -1262
rect 562 -1396 630 -1318
rect 754 -1102 822 -1070
rect 754 -1158 760 -1102
rect 816 -1158 822 -1102
rect 754 -1182 822 -1158
rect 754 -1238 760 -1182
rect 816 -1238 822 -1182
rect 754 -1262 822 -1238
rect 754 -1318 760 -1262
rect 816 -1318 822 -1262
rect 754 -1396 822 -1318
rect 946 -1102 1014 -1070
rect 946 -1158 952 -1102
rect 1008 -1158 1014 -1102
rect 946 -1182 1014 -1158
rect 946 -1238 952 -1182
rect 1008 -1238 1014 -1182
rect 946 -1262 1014 -1238
rect 946 -1318 952 -1262
rect 1008 -1318 1014 -1262
rect 946 -1396 1014 -1318
rect 1138 -1102 1206 -1070
rect 1138 -1158 1144 -1102
rect 1200 -1158 1206 -1102
rect 1138 -1182 1206 -1158
rect 1138 -1238 1144 -1182
rect 1200 -1238 1206 -1182
rect 1138 -1262 1206 -1238
rect 1138 -1318 1144 -1262
rect 1200 -1318 1206 -1262
rect 1138 -1396 1206 -1318
rect 1330 -1102 1398 -1070
rect 1330 -1158 1336 -1102
rect 1392 -1158 1398 -1102
rect 1330 -1182 1398 -1158
rect 1330 -1238 1336 -1182
rect 1392 -1238 1398 -1182
rect 1330 -1262 1398 -1238
rect 1330 -1318 1336 -1262
rect 1392 -1318 1398 -1262
rect 1330 -1396 1398 -1318
rect 1522 -1102 1590 -1070
rect 1522 -1158 1528 -1102
rect 1584 -1158 1590 -1102
rect 1522 -1182 1590 -1158
rect 1522 -1238 1528 -1182
rect 1584 -1238 1590 -1182
rect 1522 -1262 1590 -1238
rect 1522 -1318 1528 -1262
rect 1584 -1318 1590 -1262
rect 1522 -1396 1590 -1318
rect 1714 -1102 1782 -1070
rect 1714 -1158 1720 -1102
rect 1776 -1158 1782 -1102
rect 1714 -1182 1782 -1158
rect 1714 -1238 1720 -1182
rect 1776 -1238 1782 -1182
rect 1714 -1262 1782 -1238
rect 1714 -1318 1720 -1262
rect 1776 -1318 1782 -1262
rect 1714 -1396 1782 -1318
rect 1906 -1102 1974 -1072
rect 1906 -1158 1912 -1102
rect 1968 -1158 1974 -1102
rect 1906 -1182 1974 -1158
rect 1906 -1238 1912 -1182
rect 1968 -1238 1974 -1182
rect 1906 -1262 1974 -1238
rect 1906 -1318 1912 -1262
rect 1968 -1318 1974 -1262
rect 1906 -1396 1974 -1318
rect 2098 -1102 2166 -1070
rect 2098 -1158 2104 -1102
rect 2160 -1158 2166 -1102
rect 2098 -1182 2166 -1158
rect 2098 -1238 2104 -1182
rect 2160 -1238 2166 -1182
rect 2098 -1262 2166 -1238
rect 2098 -1318 2104 -1262
rect 2160 -1318 2166 -1262
rect 2098 -1396 2166 -1318
rect 2290 -1102 2358 -1070
rect 2290 -1158 2296 -1102
rect 2352 -1158 2358 -1102
rect 2290 -1182 2358 -1158
rect 2290 -1238 2296 -1182
rect 2352 -1238 2358 -1182
rect 2290 -1262 2358 -1238
rect 2290 -1318 2296 -1262
rect 2352 -1318 2358 -1262
rect 2290 -1396 2358 -1318
rect 2482 -1102 2550 -1072
rect 2482 -1158 2488 -1102
rect 2544 -1158 2550 -1102
rect 2482 -1182 2550 -1158
rect 2482 -1238 2488 -1182
rect 2544 -1238 2550 -1182
rect 2482 -1262 2550 -1238
rect 2482 -1318 2488 -1262
rect 2544 -1318 2550 -1262
rect 2482 -1396 2550 -1318
rect 2674 -1102 2742 -1070
rect 2674 -1158 2680 -1102
rect 2736 -1158 2742 -1102
rect 2674 -1182 2742 -1158
rect 2674 -1238 2680 -1182
rect 2736 -1238 2742 -1182
rect 2674 -1262 2742 -1238
rect 2674 -1318 2680 -1262
rect 2736 -1318 2742 -1262
rect 2674 -1396 2742 -1318
rect 2866 -1102 2934 -1072
rect 2866 -1158 2872 -1102
rect 2928 -1158 2934 -1102
rect 2866 -1182 2934 -1158
rect 2866 -1238 2872 -1182
rect 2928 -1238 2934 -1182
rect 2866 -1262 2934 -1238
rect 2866 -1318 2872 -1262
rect 2928 -1318 2934 -1262
rect 2866 -1396 2934 -1318
rect 3058 -1102 3126 -1070
rect 3058 -1158 3064 -1102
rect 3120 -1158 3126 -1102
rect 3058 -1182 3126 -1158
rect 3058 -1238 3064 -1182
rect 3120 -1238 3126 -1182
rect 3058 -1262 3126 -1238
rect 3058 -1318 3064 -1262
rect 3120 -1318 3126 -1262
rect 3058 -1396 3126 -1318
rect 3250 -1102 3318 -1070
rect 3250 -1158 3256 -1102
rect 3312 -1158 3318 -1102
rect 3250 -1182 3318 -1158
rect 3250 -1238 3256 -1182
rect 3312 -1238 3318 -1182
rect 3250 -1262 3318 -1238
rect 3250 -1318 3256 -1262
rect 3312 -1318 3318 -1262
rect 3250 -1396 3318 -1318
rect 3442 -1102 3510 -1070
rect 3442 -1158 3448 -1102
rect 3504 -1158 3510 -1102
rect 3442 -1182 3510 -1158
rect 3442 -1238 3448 -1182
rect 3504 -1238 3510 -1182
rect 3442 -1262 3510 -1238
rect 3442 -1318 3448 -1262
rect 3504 -1318 3510 -1262
rect 3442 -1396 3510 -1318
rect 3634 -1102 3702 -1070
rect 3634 -1158 3640 -1102
rect 3696 -1158 3702 -1102
rect 3634 -1182 3702 -1158
rect 3634 -1238 3640 -1182
rect 3696 -1238 3702 -1182
rect 3634 -1262 3702 -1238
rect 3634 -1318 3640 -1262
rect 3696 -1318 3702 -1262
rect 3634 -1396 3702 -1318
rect 3826 -1102 3894 -1070
rect 3826 -1158 3832 -1102
rect 3888 -1158 3894 -1102
rect 3826 -1182 3894 -1158
rect 3826 -1238 3832 -1182
rect 3888 -1238 3894 -1182
rect 3826 -1262 3894 -1238
rect 3826 -1318 3832 -1262
rect 3888 -1318 3894 -1262
rect 3826 -1396 3894 -1318
rect 4018 -1102 4086 -1070
rect 4018 -1158 4024 -1102
rect 4080 -1158 4086 -1102
rect 4018 -1182 4086 -1158
rect 4018 -1238 4024 -1182
rect 4080 -1238 4086 -1182
rect 4018 -1262 4086 -1238
rect 4018 -1318 4024 -1262
rect 4080 -1318 4086 -1262
rect 4018 -1396 4086 -1318
rect 178 -1450 4088 -1396
rect 78 -1640 4180 -1450
use sky130_fd_pr__pfet_01v8_CC7KEW  sky130_fd_pr__pfet_01v8_CC7KEW_0
timestamp 1627926120
transform 1 0 2131 0 1 -1038
box -2081 -400 2081 400
<< labels >>
rlabel locali s 276 -1706 2286 -1502 4 GND
rlabel metal3 s 82 -1636 4176 -1558 4 vh
port 1 nsew
rlabel metal1 s 134 -1430 4034 -1378 4 gate
port 2 nsew
rlabel metal2 s 90 -612 4174 -524 4 VDD
port 3 nsew
<< end >>
