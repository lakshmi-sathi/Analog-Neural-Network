magic
tech sky130A
magscale 1 2
timestamp 1624087956
<< error_s >>
rect 135695 581948 135730 582332
rect 135809 582046 135844 582332
rect 135927 582046 135962 582332
rect 136045 582046 136080 582332
rect 136163 582046 136198 582332
rect 136281 582046 136316 582332
rect 136399 582046 136434 582332
rect 136517 582046 136552 582332
rect 136635 582046 136670 582332
rect 136753 582046 136788 582332
rect 136871 582046 136906 582332
rect 136989 582046 137024 582332
rect 137107 582046 137142 582332
rect 137225 582046 137260 582332
rect 137343 582046 137378 582332
rect 137461 582046 137496 582332
rect 137579 582046 137614 582332
rect 137697 582046 137732 582332
rect 137815 582046 137850 582332
rect 137933 582046 137968 582332
rect 138051 582046 138086 582332
rect 138169 582046 138204 582332
rect 138287 582046 138322 582332
rect 138405 582046 138440 582332
rect 138523 582046 138558 582332
rect 138641 582046 138676 582332
rect 138759 582046 138793 582332
rect 138876 582046 138911 582332
rect 138994 582046 139029 582332
rect 139112 582046 139147 582332
rect 139230 582046 139265 582332
rect 139348 582046 139383 582332
rect 139466 582046 139501 582332
rect 139584 582046 139619 582332
rect 139702 582046 139737 582332
rect 139820 582046 139855 582332
rect 139938 582046 139973 582332
rect 140056 582046 140091 582332
rect 140174 582046 140209 582332
rect 140292 582046 140327 582332
rect 140410 582046 140445 582332
rect 140528 582046 140563 582332
rect 140646 582046 140681 582332
rect 140764 582046 140799 582332
rect 140882 582046 140917 582332
rect 141000 582046 141035 582332
rect 141118 582046 141120 582332
rect 135695 581947 135729 581948
rect 135792 581885 141120 581886
rect 135791 581851 141120 581885
rect 135791 581569 141120 581603
rect 135792 581568 141120 581569
rect 135695 581506 135729 581507
rect 135695 579898 135730 581506
rect 135809 580832 135844 581408
rect 135927 580832 135962 581408
rect 136045 580832 136080 581408
rect 136163 580832 136198 581408
rect 136281 580832 136316 581408
rect 136399 580832 136434 581408
rect 136517 580832 136552 581408
rect 136635 580832 136670 581408
rect 136753 580832 136788 581408
rect 136871 580832 136906 581408
rect 136989 580832 137024 581408
rect 137107 580832 137142 581408
rect 137225 580832 137260 581408
rect 137343 580832 137378 581408
rect 137461 580832 137496 581408
rect 137579 580832 137614 581408
rect 137697 580832 137732 581408
rect 137815 580832 137850 581408
rect 137933 580832 137968 581408
rect 138051 580832 138086 581408
rect 138169 580832 138204 581408
rect 138287 580832 138322 581408
rect 138405 580832 138440 581408
rect 138523 580832 138558 581408
rect 138641 580832 138676 581408
rect 138759 580832 138793 581408
rect 138876 580832 138911 581408
rect 138994 580832 139029 581408
rect 139112 580832 139147 581408
rect 139230 580832 139265 581408
rect 139348 580832 139383 581408
rect 139466 580832 139501 581408
rect 139584 580832 139619 581408
rect 139702 580832 139737 581408
rect 139820 580832 139855 581408
rect 139938 580832 139973 581408
rect 140056 580832 140091 581408
rect 140174 580832 140209 581408
rect 140292 580832 140327 581408
rect 140410 580832 140445 581408
rect 140528 580832 140563 581408
rect 140646 580832 140681 581408
rect 140764 580832 140799 581408
rect 140882 580832 140917 581408
rect 141000 580832 141035 581408
rect 141118 580832 141120 581408
rect 135868 580738 135902 580773
rect 135986 580738 136020 580773
rect 136104 580738 136138 580773
rect 136222 580738 136256 580773
rect 136340 580738 136374 580773
rect 136458 580738 136492 580773
rect 136576 580738 136610 580773
rect 136694 580738 136728 580773
rect 136812 580738 136846 580773
rect 136930 580738 136964 580773
rect 137048 580738 137082 580773
rect 137166 580738 137200 580773
rect 137284 580738 137318 580773
rect 137402 580738 137436 580773
rect 137520 580738 137554 580773
rect 137638 580738 137672 580773
rect 137756 580738 137790 580773
rect 137874 580738 137908 580773
rect 137992 580738 138026 580773
rect 138110 580738 138144 580773
rect 138228 580738 138262 580773
rect 138346 580738 138380 580773
rect 138464 580738 138498 580773
rect 138582 580738 138616 580773
rect 138700 580738 138734 580773
rect 138818 580738 138852 580773
rect 138936 580738 138970 580773
rect 139054 580738 139088 580773
rect 139172 580738 139206 580773
rect 139290 580738 139324 580773
rect 139408 580738 139442 580773
rect 139526 580738 139560 580773
rect 139644 580738 139678 580773
rect 139762 580738 139796 580773
rect 139880 580738 139914 580773
rect 139998 580738 140032 580773
rect 140116 580738 140150 580773
rect 140234 580738 140268 580773
rect 140352 580738 140386 580773
rect 140470 580738 140504 580773
rect 140588 580738 140622 580773
rect 140706 580738 140740 580773
rect 140824 580738 140858 580773
rect 140942 580738 140976 580773
rect 141060 580738 141094 580773
rect 135868 580631 135902 580666
rect 135986 580631 136020 580666
rect 136104 580631 136138 580666
rect 136222 580631 136256 580666
rect 136340 580631 136374 580666
rect 136458 580631 136492 580666
rect 136576 580631 136610 580666
rect 136694 580631 136728 580666
rect 136812 580631 136846 580666
rect 136930 580631 136964 580666
rect 137048 580631 137082 580666
rect 137166 580631 137200 580666
rect 137284 580631 137318 580666
rect 137402 580631 137436 580666
rect 137520 580631 137554 580666
rect 137638 580631 137672 580666
rect 137756 580631 137790 580666
rect 137874 580631 137908 580666
rect 137992 580631 138026 580666
rect 138110 580631 138144 580666
rect 138228 580631 138262 580666
rect 138346 580631 138380 580666
rect 138464 580631 138498 580666
rect 138582 580631 138616 580666
rect 138700 580631 138734 580666
rect 138818 580631 138852 580666
rect 138936 580631 138970 580666
rect 139054 580631 139088 580666
rect 139172 580631 139206 580666
rect 139290 580631 139324 580666
rect 139408 580631 139442 580666
rect 139526 580631 139560 580666
rect 139644 580631 139678 580666
rect 139762 580631 139796 580666
rect 139880 580631 139914 580666
rect 139998 580631 140032 580666
rect 140116 580631 140150 580666
rect 140234 580631 140268 580666
rect 140352 580631 140386 580666
rect 140470 580631 140504 580666
rect 140588 580631 140622 580666
rect 140706 580631 140740 580666
rect 140824 580631 140858 580666
rect 140942 580631 140976 580666
rect 141060 580631 141094 580666
rect 135809 579996 135844 580572
rect 135927 579996 135962 580572
rect 136045 579996 136080 580572
rect 136163 579996 136198 580572
rect 136281 579996 136316 580572
rect 136399 579996 136434 580572
rect 136517 579996 136552 580572
rect 136635 579996 136670 580572
rect 136753 579996 136788 580572
rect 136871 579996 136906 580572
rect 136989 579996 137024 580572
rect 137107 579996 137142 580572
rect 137225 579996 137260 580572
rect 137343 579996 137378 580572
rect 137461 579996 137496 580572
rect 137579 579996 137614 580572
rect 137697 579996 137732 580572
rect 137815 579996 137850 580572
rect 137933 579996 137968 580572
rect 138051 579996 138086 580572
rect 138169 579996 138204 580572
rect 138287 579996 138322 580572
rect 138405 579996 138440 580572
rect 138523 579996 138558 580572
rect 138641 579996 138676 580572
rect 138759 579996 138793 580572
rect 138876 579996 138911 580572
rect 138994 579996 139029 580572
rect 139112 579996 139147 580572
rect 139230 579996 139265 580572
rect 139348 579996 139383 580572
rect 139466 579996 139501 580572
rect 139584 579996 139619 580572
rect 139702 579996 139737 580572
rect 139820 579996 139855 580572
rect 139938 579996 139973 580572
rect 140056 579996 140091 580572
rect 140174 579996 140209 580572
rect 140292 579996 140327 580572
rect 140410 579996 140445 580572
rect 140528 579996 140563 580572
rect 140646 579996 140681 580572
rect 140764 579996 140799 580572
rect 140882 579996 140917 580572
rect 141000 579996 141035 580572
rect 141118 579996 141120 580572
rect 181482 580322 181488 580327
rect 183036 580322 183042 580327
rect 181476 580315 181481 580321
rect 183043 580315 183048 580321
rect 135695 579897 135729 579898
rect 135659 579589 141120 579842
rect 136753 579358 136754 579374
rect 136871 579358 136872 579374
rect 136989 579358 136990 579374
rect 137107 579358 137108 579374
rect 136045 578782 136080 579358
rect 136163 578782 136198 579358
rect 136281 578782 136316 579358
rect 136399 578782 136434 579358
rect 136517 578782 136552 579358
rect 136635 578782 136670 579358
rect 136737 579342 136788 579358
rect 136855 579342 136906 579358
rect 136973 579342 137024 579358
rect 137091 579342 137142 579358
rect 136753 578798 136788 579342
rect 136871 578798 136906 579342
rect 136989 578798 137024 579342
rect 137107 578798 137142 579342
rect 136737 578782 136788 578798
rect 136855 578782 136906 578798
rect 136973 578782 137024 578798
rect 137091 578782 137142 578798
rect 137225 578782 137260 579358
rect 137343 578782 137378 579358
rect 137461 578782 137496 579358
rect 137579 578782 137614 579358
rect 137697 578782 137732 579358
rect 137815 578782 137850 579358
rect 137933 578782 137968 579358
rect 138051 578782 138086 579358
rect 138169 578782 138204 579358
rect 138287 578782 138322 579358
rect 138405 578782 138440 579358
rect 138523 578782 138558 579358
rect 138641 578782 138676 579358
rect 138758 578782 138759 578816
rect 136753 578766 136754 578782
rect 136871 578766 136872 578782
rect 136989 578766 136990 578782
rect 137107 578766 137108 578782
rect 138792 578766 138794 579374
rect 140090 579358 140091 579374
rect 140208 579358 140209 579374
rect 140326 579358 140327 579374
rect 140444 579358 140445 579374
rect 140562 579358 140563 579374
rect 140680 579358 140681 579374
rect 140798 579358 140799 579374
rect 140916 579358 140917 579374
rect 141034 579358 141035 579374
rect 138876 578782 138911 579358
rect 138994 578782 139029 579358
rect 139112 578782 139147 579358
rect 139230 578782 139265 579358
rect 139348 578782 139383 579358
rect 139466 578782 139501 579358
rect 139584 578782 139619 579358
rect 139702 578782 139737 579358
rect 139820 578782 139855 579358
rect 139938 578782 139973 579358
rect 140056 579342 140107 579358
rect 140174 579342 140225 579358
rect 140292 579342 140343 579358
rect 140410 579342 140461 579358
rect 140528 579342 140579 579358
rect 140646 579342 140697 579358
rect 140764 579342 140815 579358
rect 140882 579342 140933 579358
rect 141000 579342 141051 579358
rect 140056 578798 140091 579342
rect 140174 578798 140209 579342
rect 140292 578798 140327 579342
rect 140410 578798 140445 579342
rect 140528 578798 140563 579342
rect 140646 578798 140681 579342
rect 140764 578798 140799 579342
rect 140882 578798 140917 579342
rect 141000 578798 141035 579342
rect 140056 578782 140107 578798
rect 140174 578782 140225 578798
rect 140292 578782 140343 578798
rect 140410 578782 140461 578798
rect 140528 578782 140579 578798
rect 140646 578782 140697 578798
rect 140764 578782 140815 578798
rect 140882 578782 140933 578798
rect 141000 578782 141051 578798
rect 141118 578782 141120 579358
rect 140090 578766 140091 578782
rect 140208 578766 140209 578782
rect 140326 578766 140327 578782
rect 140444 578766 140445 578782
rect 140562 578766 140563 578782
rect 140680 578766 140681 578782
rect 140798 578766 140799 578782
rect 140916 578766 140917 578782
rect 141034 578766 141035 578782
rect 135868 578688 135902 578723
rect 135986 578688 136020 578723
rect 136104 578688 136138 578723
rect 136222 578688 136256 578723
rect 136340 578688 136374 578723
rect 136458 578688 136492 578723
rect 136576 578688 136610 578723
rect 136694 578688 136728 578723
rect 136812 578688 136846 578723
rect 136930 578688 136964 578723
rect 137048 578688 137082 578723
rect 137166 578688 137200 578723
rect 137284 578688 137318 578723
rect 137402 578688 137436 578723
rect 137520 578688 137554 578723
rect 137638 578688 137672 578723
rect 137756 578688 137790 578723
rect 137874 578688 137908 578723
rect 137992 578688 138026 578723
rect 138110 578688 138144 578723
rect 138228 578688 138262 578723
rect 138346 578688 138380 578723
rect 138464 578688 138498 578723
rect 138582 578688 138616 578723
rect 138700 578688 138734 578723
rect 138818 578688 138852 578723
rect 138936 578688 138970 578723
rect 139054 578688 139088 578723
rect 139172 578688 139206 578723
rect 139290 578688 139324 578723
rect 139408 578688 139442 578723
rect 139526 578688 139560 578723
rect 139644 578688 139678 578723
rect 139762 578688 139796 578723
rect 139880 578688 139914 578723
rect 139998 578688 140032 578723
rect 140116 578688 140150 578723
rect 140234 578688 140268 578723
rect 140352 578688 140386 578723
rect 140470 578688 140504 578723
rect 140588 578688 140622 578723
rect 140706 578688 140740 578723
rect 140824 578688 140858 578723
rect 140942 578688 140976 578723
rect 141060 578688 141094 578723
rect 135868 578581 135902 578616
rect 135986 578581 136020 578616
rect 136104 578581 136138 578616
rect 136222 578581 136256 578616
rect 136340 578581 136374 578616
rect 136458 578581 136492 578616
rect 136576 578581 136610 578616
rect 136694 578581 136728 578616
rect 136812 578581 136846 578616
rect 136930 578581 136964 578616
rect 137048 578581 137082 578616
rect 137166 578581 137200 578616
rect 137284 578581 137318 578616
rect 137402 578581 137436 578616
rect 137520 578581 137554 578616
rect 137638 578581 137672 578616
rect 137756 578581 137790 578616
rect 137874 578581 137908 578616
rect 137992 578581 138026 578616
rect 138110 578581 138144 578616
rect 138228 578581 138262 578616
rect 138346 578581 138380 578616
rect 138464 578581 138498 578616
rect 138582 578581 138616 578616
rect 138700 578581 138734 578616
rect 138818 578581 138852 578616
rect 138936 578581 138970 578616
rect 139054 578581 139088 578616
rect 139172 578581 139206 578616
rect 139290 578581 139324 578616
rect 139408 578581 139442 578616
rect 139526 578581 139560 578616
rect 139644 578581 139678 578616
rect 139762 578581 139796 578616
rect 139880 578581 139914 578616
rect 139998 578581 140032 578616
rect 140116 578581 140150 578616
rect 140234 578581 140268 578616
rect 140352 578581 140386 578616
rect 140470 578581 140504 578616
rect 140588 578581 140622 578616
rect 140706 578581 140740 578616
rect 140824 578581 140858 578616
rect 140942 578581 140976 578616
rect 141060 578581 141094 578616
rect 136753 578522 136754 578538
rect 136871 578522 136872 578538
rect 136989 578522 136990 578538
rect 137107 578522 137108 578538
rect 135809 577946 135844 578522
rect 135927 577946 135962 578522
rect 136045 577946 136080 578522
rect 136163 577946 136198 578522
rect 136281 577946 136316 578522
rect 136399 577946 136434 578522
rect 136517 577946 136552 578522
rect 136635 577946 136670 578522
rect 136737 578506 136788 578522
rect 136855 578506 136906 578522
rect 136973 578506 137024 578522
rect 137091 578506 137142 578522
rect 136753 577962 136788 578506
rect 136871 577962 136906 578506
rect 136989 577962 137024 578506
rect 137107 577962 137142 578506
rect 136737 577946 136788 577962
rect 136855 577946 136906 577962
rect 136973 577946 137024 577962
rect 137091 577946 137142 577962
rect 137225 577946 137260 578522
rect 137343 577946 137378 578522
rect 137461 577946 137496 578522
rect 137579 577946 137614 578522
rect 137697 577946 137732 578522
rect 137815 577946 137850 578522
rect 137933 577946 137968 578522
rect 138051 577946 138086 578522
rect 138169 577946 138204 578522
rect 138287 577946 138322 578522
rect 138405 577946 138440 578522
rect 138523 577946 138558 578522
rect 138641 577946 138676 578522
rect 138758 577946 138759 577980
rect 136753 577930 136754 577946
rect 136871 577930 136872 577946
rect 136989 577930 136990 577946
rect 137107 577930 137108 577946
rect 138792 577930 138794 578538
rect 140090 578522 140091 578538
rect 140208 578522 140209 578538
rect 140326 578522 140327 578538
rect 140444 578522 140445 578538
rect 140562 578522 140563 578538
rect 140680 578522 140681 578538
rect 140798 578522 140799 578538
rect 140916 578522 140917 578538
rect 141034 578522 141035 578538
rect 138876 577946 138911 578522
rect 138994 577946 139029 578522
rect 139112 577946 139147 578522
rect 139230 577946 139265 578522
rect 139348 577946 139383 578522
rect 139466 577946 139501 578522
rect 139584 577946 139619 578522
rect 139702 577946 139737 578522
rect 139820 577946 139855 578522
rect 139938 577946 139973 578522
rect 140056 578506 140107 578522
rect 140174 578506 140225 578522
rect 140292 578506 140343 578522
rect 140410 578506 140461 578522
rect 140528 578506 140579 578522
rect 140646 578506 140697 578522
rect 140764 578506 140815 578522
rect 140882 578506 140933 578522
rect 141000 578506 141051 578522
rect 140056 577962 140091 578506
rect 140174 577962 140209 578506
rect 140292 577962 140327 578506
rect 140410 577962 140445 578506
rect 140528 577962 140563 578506
rect 140646 577962 140681 578506
rect 140764 577962 140799 578506
rect 140882 577962 140917 578506
rect 141000 577962 141035 578506
rect 140056 577946 140107 577962
rect 140174 577946 140225 577962
rect 140292 577946 140343 577962
rect 140410 577946 140461 577962
rect 140528 577946 140579 577962
rect 140646 577946 140697 577962
rect 140764 577946 140815 577962
rect 140882 577946 140933 577962
rect 141000 577946 141051 577962
rect 141118 577946 141120 578522
rect 140090 577930 140091 577946
rect 140208 577930 140209 577946
rect 140326 577930 140327 577946
rect 140444 577930 140445 577946
rect 140562 577930 140563 577946
rect 140680 577930 140681 577946
rect 140798 577930 140799 577946
rect 140916 577930 140917 577946
rect 141034 577930 141035 577946
rect 80675 577130 80691 577131
rect 80693 577130 80709 577131
rect 80823 577130 80839 577131
rect 80841 577130 80857 577131
rect 80971 577130 80987 577131
rect 80989 577130 81005 577131
rect 81119 577130 81135 577131
rect 81137 577130 81153 577131
rect 81267 577130 81283 577131
rect 81285 577130 81301 577131
rect 81415 577130 81431 577131
rect 81433 577130 81449 577131
rect 81563 577130 81579 577131
rect 81581 577130 81597 577131
rect 81711 577130 81727 577131
rect 81729 577130 81745 577131
rect 81859 577130 81875 577131
rect 81877 577130 81893 577131
rect 82007 577130 82023 577131
rect 82025 577130 82041 577131
rect 82155 577130 82171 577131
rect 82173 577130 82189 577131
rect 82303 577130 82319 577131
rect 82321 577130 82337 577131
rect 82451 577130 82467 577131
rect 82469 577130 82485 577131
rect 82599 577130 82615 577131
rect 82617 577130 82633 577131
rect 82747 577130 82763 577131
rect 82765 577130 82781 577131
rect 82895 577130 82911 577131
rect 82913 577130 82929 577131
rect 83043 577130 83059 577131
rect 83061 577130 83077 577131
rect 83191 577130 83207 577131
rect 83209 577130 83225 577131
rect 83339 577130 83355 577131
rect 83357 577130 83373 577131
rect 83487 577130 83503 577131
rect 83505 577130 83521 577131
rect 83635 577130 83651 577131
rect 83653 577130 83669 577131
rect 83783 577130 83799 577131
rect 83801 577130 83817 577131
rect 83931 577130 83947 577131
rect 83949 577130 83965 577131
rect 84079 577130 84095 577131
rect 84097 577130 84113 577131
rect 84227 577130 84243 577131
rect 84245 577130 84261 577131
rect 84375 577130 84391 577131
rect 84393 577130 84409 577131
rect 84523 577130 84539 577131
rect 84541 577130 84557 577131
rect 84671 577130 84687 577131
rect 84689 577130 84705 577131
rect 84819 577130 84835 577131
rect 84837 577130 84853 577131
rect 84967 577130 84983 577131
rect 84985 577130 85001 577131
rect 85115 577130 85131 577131
rect 85133 577130 85149 577131
rect 85263 577130 85279 577131
rect 85281 577130 85297 577131
rect 85411 577130 85427 577131
rect 85429 577130 85445 577131
rect 85559 577130 85575 577131
rect 85577 577130 85593 577131
rect 85707 577130 85723 577131
rect 85725 577130 85741 577131
rect 85855 577130 85871 577131
rect 85873 577130 85889 577131
rect 86003 577130 86019 577131
rect 86021 577130 86037 577131
rect 86151 577130 86167 577131
rect 86169 577130 86185 577131
rect 86299 577130 86315 577131
rect 86317 577130 86333 577131
rect 86447 577130 86463 577131
rect 86465 577130 86481 577131
rect 86595 577130 86611 577131
rect 86613 577130 86629 577131
rect 86743 577130 86759 577131
rect 86761 577130 86777 577131
rect 86891 577130 86907 577131
rect 86909 577130 86925 577131
rect 87039 577130 87055 577131
rect 87057 577130 87073 577131
rect 87187 577130 87203 577131
rect 87205 577130 87221 577131
rect 87335 577130 87351 577131
rect 87353 577130 87369 577131
rect 87483 577130 87499 577131
rect 87501 577130 87517 577131
rect 87631 577130 87647 577131
rect 87649 577130 87665 577131
rect 87779 577130 87795 577131
rect 87797 577130 87813 577131
rect 87927 577130 87943 577131
rect 87945 577130 87961 577131
rect 88075 577130 88091 577131
rect 88093 577130 88109 577131
rect 88223 577130 88239 577131
rect 88241 577130 88257 577131
rect 88371 577130 88387 577131
rect 88389 577130 88405 577131
rect 88519 577130 88535 577131
rect 88537 577130 88553 577131
rect 88667 577130 88683 577131
rect 88685 577130 88701 577131
rect 88815 577130 88831 577131
rect 88833 577130 88849 577131
rect 88963 577130 88979 577131
rect 88981 577130 88997 577131
rect 89111 577130 89127 577131
rect 89129 577130 89145 577131
rect 89259 577130 89275 577131
rect 89277 577130 89293 577131
rect 89407 577130 89423 577131
rect 89425 577130 89441 577131
rect 89555 577130 89571 577131
rect 89573 577130 89589 577131
rect 89703 577130 89719 577131
rect 89721 577130 89737 577131
rect 137347 577130 137363 577131
rect 137365 577130 137381 577131
rect 137465 577130 137481 577131
rect 137483 577130 137499 577131
rect 137583 577130 137599 577131
rect 137601 577130 137617 577131
rect 137701 577130 137717 577131
rect 137719 577130 137735 577131
rect 138873 577130 138889 577131
rect 138891 577130 138907 577131
rect 138991 577130 139007 577131
rect 139009 577130 139025 577131
rect 139109 577130 139125 577131
rect 139127 577130 139143 577131
rect 139227 577130 139243 577131
rect 139245 577130 139261 577131
rect 139345 577130 139361 577131
rect 139363 577130 139379 577131
rect 139463 577130 139479 577131
rect 139481 577130 139497 577131
rect 139581 577130 139597 577131
rect 139599 577130 139615 577131
rect 139699 577130 139715 577131
rect 139717 577130 139733 577131
rect 139817 577130 139833 577131
rect 139835 577130 139851 577131
rect 139935 577130 139951 577131
rect 139953 577130 139969 577131
rect 140053 577130 140069 577131
rect 140071 577130 140087 577131
rect 140171 577130 140187 577131
rect 140189 577130 140205 577131
rect 140289 577130 140305 577131
rect 140307 577130 140323 577131
rect 140407 577130 140423 577131
rect 140425 577130 140441 577131
rect 140525 577130 140541 577131
rect 140543 577130 140559 577131
rect 140643 577130 140659 577131
rect 140661 577130 140677 577131
rect 144717 577130 144733 577131
rect 144735 577130 144751 577131
rect 144865 577130 144881 577131
rect 144883 577130 144899 577131
rect 145013 577130 145029 577131
rect 145031 577130 145047 577131
rect 145161 577130 145177 577131
rect 145179 577130 145195 577131
rect 145309 577130 145325 577131
rect 145327 577130 145343 577131
rect 145457 577130 145473 577131
rect 145475 577130 145491 577131
rect 145605 577130 145621 577131
rect 145623 577130 145639 577131
rect 145753 577130 145769 577131
rect 145771 577130 145787 577131
rect 80675 577115 80676 577130
rect 80823 577115 80824 577130
rect 80971 577115 80972 577130
rect 81119 577115 81120 577130
rect 81267 577115 81268 577130
rect 81415 577115 81416 577130
rect 81563 577115 81564 577130
rect 81711 577115 81712 577130
rect 81859 577115 81860 577130
rect 82007 577115 82008 577130
rect 82155 577115 82156 577130
rect 82303 577115 82304 577130
rect 82451 577115 82452 577130
rect 82599 577115 82600 577130
rect 82747 577115 82748 577130
rect 82895 577115 82896 577130
rect 83043 577115 83044 577130
rect 83191 577115 83192 577130
rect 83339 577115 83340 577130
rect 83487 577115 83488 577130
rect 83635 577115 83636 577130
rect 83783 577115 83784 577130
rect 83931 577115 83932 577130
rect 84079 577115 84080 577130
rect 84227 577115 84228 577130
rect 84375 577115 84376 577130
rect 84523 577115 84524 577130
rect 84671 577115 84672 577130
rect 84852 577115 84853 577130
rect 85000 577115 85001 577130
rect 85148 577115 85149 577130
rect 85296 577115 85297 577130
rect 85444 577115 85445 577130
rect 85592 577115 85593 577130
rect 85740 577115 85741 577130
rect 85888 577115 85889 577130
rect 86036 577115 86037 577130
rect 86184 577115 86185 577130
rect 86332 577115 86333 577130
rect 86480 577115 86481 577130
rect 86628 577115 86629 577130
rect 86776 577115 86777 577130
rect 86924 577115 86925 577130
rect 87072 577115 87073 577130
rect 87220 577115 87221 577130
rect 87368 577115 87369 577130
rect 87516 577115 87517 577130
rect 87664 577115 87665 577130
rect 87812 577115 87813 577130
rect 87960 577115 87961 577130
rect 88108 577115 88109 577130
rect 88256 577115 88257 577130
rect 88404 577115 88405 577130
rect 88552 577115 88553 577130
rect 88700 577115 88701 577130
rect 88848 577115 88849 577130
rect 88996 577115 88997 577130
rect 89144 577115 89145 577130
rect 89292 577115 89293 577130
rect 89440 577115 89441 577130
rect 89588 577115 89589 577130
rect 89736 577115 89737 577130
rect 144717 577115 144718 577130
rect 144865 577115 144866 577130
rect 145013 577115 145014 577130
rect 145161 577115 145162 577130
rect 145309 577115 145310 577130
rect 145457 577115 145458 577130
rect 145605 577115 145606 577130
rect 145753 577115 145754 577130
rect 145778 577115 145788 577130
rect 80659 577114 80709 577115
rect 80710 577114 80725 577115
rect 80659 577099 80725 577114
rect 80807 577114 80857 577115
rect 80858 577114 80873 577115
rect 80807 577099 80873 577114
rect 80955 577114 81005 577115
rect 81006 577114 81021 577115
rect 80955 577099 81021 577114
rect 81103 577114 81153 577115
rect 81154 577114 81169 577115
rect 81103 577099 81169 577114
rect 81251 577114 81301 577115
rect 81302 577114 81317 577115
rect 81251 577099 81317 577114
rect 81399 577114 81449 577115
rect 81450 577114 81465 577115
rect 81399 577099 81465 577114
rect 81547 577114 81597 577115
rect 81598 577114 81613 577115
rect 81547 577099 81613 577114
rect 81695 577114 81745 577115
rect 81746 577114 81761 577115
rect 81695 577099 81761 577114
rect 81843 577114 81893 577115
rect 81894 577114 81909 577115
rect 81843 577099 81909 577114
rect 81991 577114 82041 577115
rect 82042 577114 82057 577115
rect 81991 577099 82057 577114
rect 82139 577114 82189 577115
rect 82190 577114 82205 577115
rect 82139 577099 82205 577114
rect 82287 577114 82337 577115
rect 82338 577114 82353 577115
rect 82287 577099 82353 577114
rect 82435 577114 82485 577115
rect 82486 577114 82501 577115
rect 82435 577099 82501 577114
rect 82583 577114 82633 577115
rect 82634 577114 82649 577115
rect 82583 577099 82649 577114
rect 82731 577114 82781 577115
rect 82782 577114 82797 577115
rect 82731 577099 82797 577114
rect 82879 577114 82929 577115
rect 82930 577114 82945 577115
rect 82879 577099 82945 577114
rect 83027 577114 83077 577115
rect 83078 577114 83093 577115
rect 83027 577099 83093 577114
rect 83175 577114 83225 577115
rect 83226 577114 83241 577115
rect 83175 577099 83241 577114
rect 83323 577114 83373 577115
rect 83374 577114 83389 577115
rect 83323 577099 83389 577114
rect 83471 577114 83521 577115
rect 83522 577114 83537 577115
rect 83471 577099 83537 577114
rect 83619 577114 83669 577115
rect 83670 577114 83685 577115
rect 83619 577099 83685 577114
rect 83767 577114 83817 577115
rect 83818 577114 83833 577115
rect 83767 577099 83833 577114
rect 83915 577114 83965 577115
rect 83966 577114 83981 577115
rect 83915 577099 83981 577114
rect 84063 577114 84113 577115
rect 84114 577114 84129 577115
rect 84063 577099 84129 577114
rect 84211 577114 84261 577115
rect 84262 577114 84277 577115
rect 84211 577099 84277 577114
rect 84359 577114 84409 577115
rect 84410 577114 84425 577115
rect 84359 577099 84425 577114
rect 84507 577114 84557 577115
rect 84558 577114 84573 577115
rect 84507 577099 84573 577114
rect 84655 577114 84705 577115
rect 84706 577114 84721 577115
rect 84655 577099 84721 577114
rect 84803 577114 84818 577115
rect 84819 577114 84869 577115
rect 84803 577099 84869 577114
rect 84951 577114 84966 577115
rect 84967 577114 85017 577115
rect 84951 577099 85017 577114
rect 85099 577114 85114 577115
rect 85115 577114 85165 577115
rect 85099 577099 85165 577114
rect 85247 577114 85262 577115
rect 85263 577114 85313 577115
rect 85247 577099 85313 577114
rect 85395 577114 85410 577115
rect 85411 577114 85461 577115
rect 85395 577099 85461 577114
rect 85543 577114 85558 577115
rect 85559 577114 85609 577115
rect 85543 577099 85609 577114
rect 85691 577114 85706 577115
rect 85707 577114 85757 577115
rect 85691 577099 85757 577114
rect 85839 577114 85854 577115
rect 85855 577114 85905 577115
rect 85839 577099 85905 577114
rect 85987 577114 86002 577115
rect 86003 577114 86053 577115
rect 85987 577099 86053 577114
rect 86135 577114 86150 577115
rect 86151 577114 86201 577115
rect 86135 577099 86201 577114
rect 86283 577114 86298 577115
rect 86299 577114 86349 577115
rect 86283 577099 86349 577114
rect 86431 577114 86446 577115
rect 86447 577114 86497 577115
rect 86431 577099 86497 577114
rect 86579 577114 86594 577115
rect 86595 577114 86645 577115
rect 86579 577099 86645 577114
rect 86727 577114 86742 577115
rect 86743 577114 86793 577115
rect 86727 577099 86793 577114
rect 86875 577114 86890 577115
rect 86891 577114 86941 577115
rect 86875 577099 86941 577114
rect 87023 577114 87038 577115
rect 87039 577114 87089 577115
rect 87023 577099 87089 577114
rect 87171 577114 87186 577115
rect 87187 577114 87237 577115
rect 87171 577099 87237 577114
rect 87319 577114 87334 577115
rect 87335 577114 87385 577115
rect 87319 577099 87385 577114
rect 87467 577114 87482 577115
rect 87483 577114 87533 577115
rect 87467 577099 87533 577114
rect 87615 577114 87630 577115
rect 87631 577114 87681 577115
rect 87615 577099 87681 577114
rect 87763 577114 87778 577115
rect 87779 577114 87829 577115
rect 87763 577099 87829 577114
rect 87911 577114 87926 577115
rect 87927 577114 87977 577115
rect 87911 577099 87977 577114
rect 88059 577114 88074 577115
rect 88075 577114 88125 577115
rect 88059 577099 88125 577114
rect 88207 577114 88222 577115
rect 88223 577114 88273 577115
rect 88207 577099 88273 577114
rect 88355 577114 88370 577115
rect 88371 577114 88421 577115
rect 88355 577099 88421 577114
rect 88503 577114 88518 577115
rect 88519 577114 88569 577115
rect 88503 577099 88569 577114
rect 88651 577114 88666 577115
rect 88667 577114 88717 577115
rect 88651 577099 88717 577114
rect 88799 577114 88814 577115
rect 88815 577114 88865 577115
rect 88799 577099 88865 577114
rect 88947 577114 88962 577115
rect 88963 577114 89013 577115
rect 88947 577099 89013 577114
rect 89095 577114 89110 577115
rect 89111 577114 89161 577115
rect 89095 577099 89161 577114
rect 89243 577114 89258 577115
rect 89259 577114 89309 577115
rect 89243 577099 89309 577114
rect 89391 577114 89406 577115
rect 89407 577114 89457 577115
rect 89391 577099 89457 577114
rect 89539 577114 89554 577115
rect 89555 577114 89605 577115
rect 89539 577099 89605 577114
rect 89687 577114 89702 577115
rect 89703 577114 89753 577115
rect 89687 577099 89753 577114
rect 80675 576255 80710 577099
rect 80823 576255 80858 577099
rect 80971 576255 81006 577099
rect 81119 576255 81154 577099
rect 81267 576255 81302 577099
rect 81415 576255 81450 577099
rect 81563 576255 81598 577099
rect 81711 576255 81746 577099
rect 81859 576255 81894 577099
rect 82007 576255 82042 577099
rect 82155 576255 82190 577099
rect 82303 576255 82338 577099
rect 82451 576255 82486 577099
rect 82599 576255 82634 577099
rect 82747 576255 82782 577099
rect 82895 576255 82930 577099
rect 83043 576255 83078 577099
rect 83191 576255 83226 577099
rect 83339 576255 83374 577099
rect 83487 576255 83522 577099
rect 83635 576255 83670 577099
rect 83783 576255 83818 577099
rect 83931 576255 83966 577099
rect 84079 576255 84114 577099
rect 84227 576255 84262 577099
rect 84375 576255 84410 577099
rect 84523 576255 84558 577099
rect 84671 576255 84706 577099
rect 80659 576239 80710 576255
rect 80807 576239 80858 576255
rect 80955 576239 81006 576255
rect 81103 576239 81154 576255
rect 81251 576239 81302 576255
rect 81399 576239 81450 576255
rect 81547 576239 81598 576255
rect 81695 576239 81746 576255
rect 81843 576239 81894 576255
rect 81991 576239 82042 576255
rect 82139 576239 82190 576255
rect 82287 576239 82338 576255
rect 82435 576239 82486 576255
rect 82583 576239 82634 576255
rect 82731 576239 82782 576255
rect 82879 576239 82930 576255
rect 83027 576239 83078 576255
rect 83175 576239 83226 576255
rect 83323 576239 83374 576255
rect 83471 576239 83522 576255
rect 83619 576239 83670 576255
rect 83767 576239 83818 576255
rect 83915 576239 83966 576255
rect 84063 576239 84114 576255
rect 84211 576239 84262 576255
rect 84359 576239 84410 576255
rect 84507 576239 84558 576255
rect 84655 576239 84706 576255
rect 80675 576238 80710 576239
rect 80823 576238 80858 576239
rect 80971 576238 81006 576239
rect 81119 576238 81154 576239
rect 81267 576238 81302 576239
rect 81415 576238 81450 576239
rect 81563 576238 81598 576239
rect 81711 576238 81746 576239
rect 81859 576238 81894 576239
rect 82007 576238 82042 576239
rect 82155 576238 82190 576239
rect 82303 576238 82338 576239
rect 82451 576238 82486 576239
rect 82599 576238 82634 576239
rect 82747 576238 82782 576239
rect 82895 576238 82930 576239
rect 83043 576238 83078 576239
rect 83191 576238 83226 576239
rect 83339 576238 83374 576239
rect 83487 576238 83522 576239
rect 83635 576238 83670 576239
rect 83783 576238 83818 576239
rect 83931 576238 83966 576239
rect 84079 576238 84114 576239
rect 84227 576238 84262 576239
rect 84375 576238 84410 576239
rect 84523 576238 84558 576239
rect 84671 576238 84706 576239
rect 84818 576255 84853 577099
rect 84966 576255 85001 577099
rect 85114 576255 85149 577099
rect 85262 576255 85297 577099
rect 85410 576255 85445 577099
rect 85558 576255 85593 577099
rect 85706 576255 85741 577099
rect 85854 576255 85889 577099
rect 86002 576255 86037 577099
rect 86150 576255 86185 577099
rect 86298 576255 86333 577099
rect 86446 576255 86481 577099
rect 86594 576255 86629 577099
rect 86742 576255 86777 577099
rect 86890 576255 86925 577099
rect 87038 576255 87073 577099
rect 87186 576255 87221 577099
rect 87334 576255 87369 577099
rect 87482 576255 87517 577099
rect 87630 576255 87665 577099
rect 87778 576255 87813 577099
rect 87926 576255 87961 577099
rect 88074 576255 88109 577099
rect 88222 576255 88257 577099
rect 88370 576255 88405 577099
rect 88518 576255 88553 577099
rect 88666 576255 88701 577099
rect 88814 576255 88849 577099
rect 88962 576255 88997 577099
rect 89110 576255 89145 577099
rect 89258 576255 89293 577099
rect 89406 576255 89441 577099
rect 89554 576255 89589 577099
rect 89702 576255 89737 577099
rect 84818 576239 84869 576255
rect 84966 576239 85017 576255
rect 85114 576239 85165 576255
rect 85262 576239 85313 576255
rect 85410 576239 85461 576255
rect 85558 576239 85609 576255
rect 85706 576239 85757 576255
rect 85854 576239 85905 576255
rect 86002 576239 86053 576255
rect 86150 576239 86201 576255
rect 86298 576239 86349 576255
rect 86446 576239 86497 576255
rect 86594 576239 86645 576255
rect 86742 576239 86793 576255
rect 86890 576239 86941 576255
rect 87038 576239 87089 576255
rect 87186 576239 87237 576255
rect 87334 576239 87385 576255
rect 87482 576239 87533 576255
rect 87630 576239 87681 576255
rect 87778 576239 87829 576255
rect 87926 576239 87977 576255
rect 88074 576239 88125 576255
rect 88222 576239 88273 576255
rect 88370 576239 88421 576255
rect 88518 576239 88569 576255
rect 88666 576239 88717 576255
rect 88814 576239 88865 576255
rect 88962 576239 89013 576255
rect 89110 576239 89161 576255
rect 89258 576239 89309 576255
rect 89406 576239 89457 576255
rect 89554 576239 89605 576255
rect 89702 576239 89753 576255
rect 89850 576239 89885 577114
rect 89998 576239 90033 577114
rect 90294 576239 90329 577114
rect 137111 576538 137145 577114
rect 137229 576538 137263 577114
rect 137331 577099 137397 577115
rect 137449 577099 137515 577115
rect 137567 577099 137633 577115
rect 137685 577099 137751 577115
rect 137347 576538 137381 577099
rect 137465 576538 137499 577099
rect 137583 576538 137617 577099
rect 137701 576538 137735 577099
rect 137819 576538 137853 577114
rect 137937 576538 137971 577114
rect 138055 576538 138089 577114
rect 138173 576538 138207 577114
rect 138291 576538 138325 577114
rect 138409 576538 138443 577114
rect 138527 576538 138561 577114
rect 138645 576538 138679 577114
rect 138857 577099 138923 577115
rect 138975 577099 139041 577115
rect 139093 577099 139159 577115
rect 139211 577099 139277 577115
rect 139329 577099 139395 577115
rect 139447 577099 139513 577115
rect 139565 577099 139631 577115
rect 139683 577099 139749 577115
rect 139801 577099 139867 577115
rect 139919 577099 139985 577115
rect 140037 577099 140103 577115
rect 140155 577099 140221 577115
rect 140273 577099 140339 577115
rect 140391 577099 140457 577115
rect 140509 577099 140575 577115
rect 140627 577099 140693 577115
rect 144701 577114 144751 577115
rect 144752 577114 144767 577115
rect 138873 576538 138907 577099
rect 138991 576538 139025 577099
rect 139109 576538 139143 577099
rect 139227 576538 139261 577099
rect 139345 576538 139379 577099
rect 139463 576538 139497 577099
rect 139581 576538 139615 577099
rect 139699 576538 139733 577099
rect 139817 576538 139851 577099
rect 139935 576538 139969 577099
rect 140053 576538 140087 577099
rect 140171 576538 140205 577099
rect 140289 576538 140323 577099
rect 140407 576538 140441 577099
rect 140525 576538 140559 577099
rect 140643 576538 140677 577099
rect 143316 577042 143350 577043
rect 143315 576738 143350 577042
rect 143316 576737 143350 576738
rect 143349 576681 143350 576709
rect 143349 576647 143352 576675
rect 136921 576526 136981 576527
rect 137039 576526 137099 576527
rect 137157 576526 137217 576527
rect 137275 576526 137335 576527
rect 137393 576526 137453 576527
rect 137511 576526 137571 576527
rect 137629 576526 137689 576527
rect 137747 576526 137807 576527
rect 137865 576526 137925 576527
rect 137983 576526 138043 576527
rect 138101 576526 138161 576527
rect 138219 576526 138279 576527
rect 138337 576526 138397 576527
rect 138455 576526 138515 576527
rect 138573 576526 138633 576527
rect 136934 576488 136968 576489
rect 137052 576488 137086 576489
rect 137170 576488 137204 576489
rect 137288 576488 137322 576489
rect 137406 576488 137440 576489
rect 137524 576488 137558 576489
rect 137642 576488 137676 576489
rect 136934 576455 136969 576488
rect 137052 576455 137087 576488
rect 137170 576455 137205 576488
rect 137288 576455 137323 576488
rect 137406 576455 137441 576488
rect 137524 576455 137559 576488
rect 137642 576455 137677 576488
rect 137759 576455 137795 576489
rect 137878 576488 137912 576489
rect 137996 576488 138030 576489
rect 138114 576488 138148 576489
rect 138232 576488 138266 576489
rect 138350 576488 138384 576489
rect 138468 576488 138502 576489
rect 138586 576488 138620 576489
rect 136935 576454 136969 576455
rect 137053 576454 137087 576455
rect 137171 576454 137205 576455
rect 137289 576454 137323 576455
rect 137407 576454 137441 576455
rect 137525 576454 137559 576455
rect 137643 576454 137677 576455
rect 137761 576454 137795 576455
rect 137877 576455 137912 576488
rect 137995 576455 138030 576488
rect 138113 576455 138148 576488
rect 138231 576455 138266 576488
rect 138349 576455 138384 576488
rect 138467 576455 138502 576488
rect 138585 576455 138620 576488
rect 138932 576455 138967 576488
rect 139050 576455 139085 576488
rect 139168 576455 139203 576488
rect 139286 576455 139321 576488
rect 139404 576455 139439 576488
rect 139522 576455 139557 576488
rect 139640 576455 139675 576488
rect 139757 576455 139758 576489
rect 139792 576488 139793 576489
rect 137877 576454 137911 576455
rect 137995 576454 138029 576455
rect 138113 576454 138147 576455
rect 138231 576454 138265 576455
rect 138349 576454 138383 576455
rect 138467 576454 138501 576455
rect 138585 576454 138619 576455
rect 138933 576454 138967 576455
rect 139051 576454 139085 576455
rect 139169 576454 139203 576455
rect 139287 576454 139321 576455
rect 139405 576454 139439 576455
rect 139523 576454 139557 576455
rect 139641 576454 139675 576455
rect 139759 576454 139793 576488
rect 139875 576455 139910 576488
rect 139993 576455 140028 576488
rect 140111 576455 140146 576488
rect 140229 576455 140264 576488
rect 140347 576455 140382 576488
rect 140465 576455 140500 576488
rect 140583 576455 140618 576488
rect 139875 576454 139909 576455
rect 139993 576454 140027 576455
rect 140111 576454 140145 576455
rect 140229 576454 140263 576455
rect 140347 576454 140381 576455
rect 140465 576454 140499 576455
rect 140583 576454 140617 576455
rect 136984 576438 136985 576440
rect 137102 576438 137103 576440
rect 137220 576438 137221 576440
rect 137338 576438 137339 576440
rect 137456 576438 137457 576440
rect 137574 576438 137575 576440
rect 137692 576438 137693 576440
rect 137861 576438 137862 576440
rect 137979 576438 137980 576440
rect 138097 576438 138098 576440
rect 138215 576438 138216 576440
rect 138333 576438 138334 576440
rect 138451 576438 138452 576440
rect 138569 576438 138570 576440
rect 138982 576438 138983 576440
rect 139100 576438 139101 576440
rect 139218 576438 139219 576440
rect 139336 576438 139337 576440
rect 139454 576438 139455 576440
rect 139572 576438 139573 576440
rect 139690 576438 139691 576440
rect 139859 576438 139860 576440
rect 139977 576438 139978 576440
rect 140095 576438 140096 576440
rect 140213 576438 140214 576440
rect 140331 576438 140332 576440
rect 140449 576438 140450 576440
rect 140567 576438 140568 576440
rect 136935 576381 136969 576382
rect 137053 576381 137087 576382
rect 137171 576381 137205 576382
rect 137289 576381 137323 576382
rect 137407 576381 137441 576382
rect 137525 576381 137559 576382
rect 137643 576381 137677 576382
rect 137761 576381 137795 576382
rect 137877 576381 137911 576382
rect 137995 576381 138029 576382
rect 138113 576381 138147 576382
rect 138231 576381 138265 576382
rect 138349 576381 138383 576382
rect 138467 576381 138501 576382
rect 138585 576381 138619 576382
rect 138933 576381 138967 576382
rect 139051 576381 139085 576382
rect 139169 576381 139203 576382
rect 139287 576381 139321 576382
rect 139405 576381 139439 576382
rect 139523 576381 139557 576382
rect 139641 576381 139675 576382
rect 136934 576348 136969 576381
rect 137052 576348 137087 576381
rect 137170 576348 137205 576381
rect 137288 576348 137323 576381
rect 137406 576348 137441 576381
rect 137524 576348 137559 576381
rect 137642 576348 137677 576381
rect 136934 576347 136968 576348
rect 137052 576347 137086 576348
rect 137170 576347 137204 576348
rect 137288 576347 137322 576348
rect 137406 576347 137440 576348
rect 137524 576347 137558 576348
rect 137642 576347 137676 576348
rect 137760 576347 137794 576381
rect 137877 576348 137912 576381
rect 137995 576348 138030 576381
rect 138113 576348 138148 576381
rect 138231 576348 138266 576381
rect 138349 576348 138384 576381
rect 138467 576348 138502 576381
rect 138585 576348 138620 576381
rect 138932 576348 138967 576381
rect 139050 576348 139085 576381
rect 139168 576348 139203 576381
rect 139286 576348 139321 576381
rect 139404 576348 139439 576381
rect 139522 576348 139557 576381
rect 139640 576348 139675 576381
rect 139759 576348 139793 576382
rect 139875 576381 139909 576382
rect 139993 576381 140027 576382
rect 140111 576381 140145 576382
rect 140229 576381 140263 576382
rect 140347 576381 140381 576382
rect 140465 576381 140499 576382
rect 140583 576381 140617 576382
rect 139875 576348 139910 576381
rect 139993 576348 140028 576381
rect 140111 576348 140146 576381
rect 140229 576348 140264 576381
rect 140347 576348 140382 576381
rect 140465 576348 140500 576381
rect 140583 576348 140618 576381
rect 137878 576347 137912 576348
rect 137996 576347 138030 576348
rect 138114 576347 138148 576348
rect 138232 576347 138266 576348
rect 138350 576347 138384 576348
rect 138468 576347 138502 576348
rect 138586 576347 138620 576348
rect 84818 576238 84853 576239
rect 84966 576238 85001 576239
rect 85114 576238 85149 576239
rect 85262 576238 85297 576239
rect 85410 576238 85445 576239
rect 85558 576238 85593 576239
rect 85706 576238 85741 576239
rect 85854 576238 85889 576239
rect 86002 576238 86037 576239
rect 86150 576238 86185 576239
rect 86298 576238 86333 576239
rect 86446 576238 86481 576239
rect 86594 576238 86629 576239
rect 86742 576238 86777 576239
rect 86890 576238 86925 576239
rect 87038 576238 87073 576239
rect 87186 576238 87221 576239
rect 87334 576238 87369 576239
rect 87482 576238 87517 576239
rect 87630 576238 87665 576239
rect 87778 576238 87813 576239
rect 87926 576238 87961 576239
rect 88074 576238 88109 576239
rect 88222 576238 88257 576239
rect 88370 576238 88405 576239
rect 88518 576238 88553 576239
rect 88666 576238 88701 576239
rect 88814 576238 88849 576239
rect 88962 576238 88997 576239
rect 89110 576238 89145 576239
rect 89258 576238 89293 576239
rect 89406 576238 89441 576239
rect 89554 576238 89589 576239
rect 89702 576238 89737 576239
rect 89850 576238 89884 576239
rect 89998 576238 90032 576239
rect 90294 576238 90328 576239
rect 80640 576226 80664 576227
rect 80675 576223 80676 576238
rect 80823 576223 80824 576238
rect 80971 576223 80972 576238
rect 81119 576223 81120 576238
rect 81267 576223 81268 576238
rect 81415 576223 81416 576238
rect 81563 576223 81564 576238
rect 81711 576223 81712 576238
rect 81859 576223 81860 576238
rect 82007 576223 82008 576238
rect 82155 576223 82156 576238
rect 82202 576226 82292 576227
rect 82303 576223 82304 576238
rect 82350 576226 82440 576227
rect 82451 576223 82452 576238
rect 82498 576226 82588 576227
rect 82599 576223 82600 576238
rect 82646 576226 82736 576227
rect 82747 576223 82748 576238
rect 82794 576226 82884 576227
rect 82895 576223 82896 576238
rect 82942 576226 83032 576227
rect 83043 576223 83044 576238
rect 83090 576226 83180 576227
rect 83191 576223 83192 576238
rect 83238 576226 83328 576227
rect 83339 576223 83340 576238
rect 83386 576226 83476 576227
rect 83487 576223 83488 576238
rect 83534 576226 83624 576227
rect 83635 576223 83636 576238
rect 83682 576226 83772 576227
rect 83783 576223 83784 576238
rect 83830 576226 83920 576227
rect 83931 576223 83932 576238
rect 83978 576226 84068 576227
rect 84079 576223 84080 576238
rect 84126 576226 84216 576227
rect 84227 576223 84228 576238
rect 84274 576226 84364 576227
rect 84375 576223 84376 576238
rect 84422 576226 84512 576227
rect 84523 576223 84524 576238
rect 84570 576226 84660 576227
rect 84671 576223 84672 576238
rect 84718 576226 84806 576227
rect 84852 576223 84853 576238
rect 84864 576226 84954 576227
rect 85000 576223 85001 576238
rect 85012 576226 85102 576227
rect 85148 576223 85149 576238
rect 85296 576223 85297 576238
rect 85444 576223 85445 576238
rect 85592 576223 85593 576238
rect 85740 576223 85741 576238
rect 85888 576223 85889 576238
rect 86036 576223 86037 576238
rect 86184 576223 86185 576238
rect 86332 576223 86333 576238
rect 86480 576223 86481 576238
rect 86628 576223 86629 576238
rect 86776 576223 86777 576238
rect 86924 576223 86925 576238
rect 87072 576223 87073 576238
rect 87220 576223 87221 576238
rect 87368 576223 87369 576238
rect 87516 576223 87517 576238
rect 87664 576223 87665 576238
rect 87812 576223 87813 576238
rect 87960 576223 87961 576238
rect 88108 576223 88109 576238
rect 88256 576223 88257 576238
rect 88404 576223 88405 576238
rect 88552 576223 88553 576238
rect 88700 576223 88701 576238
rect 88848 576223 88849 576238
rect 88996 576223 88997 576238
rect 89144 576223 89145 576238
rect 89292 576223 89293 576238
rect 89440 576223 89441 576238
rect 89588 576223 89589 576238
rect 89736 576223 89737 576238
rect 80640 576188 80647 576189
rect 82217 576188 82275 576189
rect 82365 576188 82423 576189
rect 82513 576188 82571 576189
rect 82661 576188 82719 576189
rect 82809 576188 82867 576189
rect 82957 576188 83015 576189
rect 83105 576188 83163 576189
rect 83253 576188 83311 576189
rect 83401 576188 83459 576189
rect 83549 576188 83607 576189
rect 83697 576188 83755 576189
rect 83845 576188 83903 576189
rect 83993 576188 84051 576189
rect 84141 576188 84199 576189
rect 84289 576188 84347 576189
rect 84437 576188 84495 576189
rect 84585 576188 84643 576189
rect 80640 576154 80648 576188
rect 80737 576155 80796 576188
rect 80885 576155 80944 576188
rect 81033 576155 81092 576188
rect 81181 576155 81240 576188
rect 81329 576155 81388 576188
rect 81477 576155 81536 576188
rect 81625 576155 81684 576188
rect 81773 576155 81832 576188
rect 81921 576155 81980 576188
rect 82069 576155 82128 576188
rect 82217 576155 82276 576188
rect 82365 576155 82424 576188
rect 82513 576155 82572 576188
rect 82661 576155 82720 576188
rect 82809 576155 82868 576188
rect 82957 576155 83016 576188
rect 83105 576155 83164 576188
rect 83253 576155 83312 576188
rect 83401 576155 83460 576188
rect 83549 576155 83608 576188
rect 83697 576155 83756 576188
rect 83845 576155 83904 576188
rect 83993 576155 84052 576188
rect 84141 576155 84200 576188
rect 84289 576155 84348 576188
rect 84437 576155 84496 576188
rect 84585 576155 84644 576188
rect 84733 576155 84791 576189
rect 84881 576188 84939 576189
rect 85029 576188 85087 576189
rect 84880 576155 84939 576188
rect 85028 576155 85087 576188
rect 85176 576155 85235 576188
rect 85324 576155 85383 576188
rect 85472 576155 85531 576188
rect 85620 576155 85679 576188
rect 85768 576155 85827 576188
rect 85916 576155 85975 576188
rect 86064 576155 86123 576188
rect 86212 576155 86271 576188
rect 86360 576155 86419 576188
rect 86508 576155 86567 576188
rect 86656 576155 86715 576188
rect 86804 576155 86863 576188
rect 86952 576155 87011 576188
rect 87100 576155 87159 576188
rect 87248 576155 87307 576188
rect 87396 576155 87455 576188
rect 87544 576155 87603 576188
rect 87692 576155 87751 576188
rect 87840 576155 87899 576188
rect 87988 576155 88047 576188
rect 88136 576155 88195 576188
rect 88284 576155 88343 576188
rect 88432 576155 88491 576188
rect 88580 576155 88639 576188
rect 88728 576155 88787 576188
rect 88876 576155 88935 576188
rect 89024 576155 89083 576188
rect 89172 576155 89231 576188
rect 89320 576155 89379 576188
rect 89468 576155 89527 576188
rect 89616 576155 89675 576188
rect 89764 576155 89823 576188
rect 89912 576155 89971 576188
rect 90060 576155 90119 576188
rect 90208 576155 90267 576188
rect 80738 576154 80796 576155
rect 80886 576154 80944 576155
rect 81034 576154 81092 576155
rect 81182 576154 81240 576155
rect 81330 576154 81388 576155
rect 81478 576154 81536 576155
rect 81626 576154 81684 576155
rect 81774 576154 81832 576155
rect 81922 576154 81980 576155
rect 82070 576154 82128 576155
rect 82218 576154 82276 576155
rect 82366 576154 82424 576155
rect 82514 576154 82572 576155
rect 82662 576154 82720 576155
rect 82810 576154 82868 576155
rect 82958 576154 83016 576155
rect 83106 576154 83164 576155
rect 83254 576154 83312 576155
rect 83402 576154 83460 576155
rect 83550 576154 83608 576155
rect 83698 576154 83756 576155
rect 83846 576154 83904 576155
rect 83994 576154 84052 576155
rect 84142 576154 84200 576155
rect 84290 576154 84348 576155
rect 84438 576154 84496 576155
rect 84586 576154 84644 576155
rect 84734 576154 84790 576155
rect 84880 576154 84938 576155
rect 85028 576154 85086 576155
rect 85176 576154 85234 576155
rect 85324 576154 85382 576155
rect 85472 576154 85530 576155
rect 85620 576154 85678 576155
rect 85768 576154 85826 576155
rect 85916 576154 85974 576155
rect 86064 576154 86122 576155
rect 86212 576154 86270 576155
rect 86360 576154 86418 576155
rect 86508 576154 86566 576155
rect 86656 576154 86714 576155
rect 86804 576154 86862 576155
rect 86952 576154 87010 576155
rect 87100 576154 87158 576155
rect 87248 576154 87306 576155
rect 87396 576154 87454 576155
rect 87544 576154 87602 576155
rect 87692 576154 87750 576155
rect 87840 576154 87898 576155
rect 87988 576154 88046 576155
rect 88136 576154 88194 576155
rect 88284 576154 88342 576155
rect 88432 576154 88490 576155
rect 88580 576154 88638 576155
rect 88728 576154 88786 576155
rect 88876 576154 88934 576155
rect 89024 576154 89082 576155
rect 89172 576154 89230 576155
rect 89320 576154 89378 576155
rect 89468 576154 89526 576155
rect 89616 576154 89674 576155
rect 89764 576154 89822 576155
rect 89912 576154 89970 576155
rect 90060 576154 90118 576155
rect 90208 576154 90266 576155
rect 80663 576138 80664 576140
rect 80811 576138 80812 576140
rect 80959 576138 80960 576140
rect 81107 576138 81108 576140
rect 81255 576138 81256 576140
rect 81403 576138 81404 576140
rect 81551 576138 81552 576140
rect 81699 576138 81700 576140
rect 81847 576138 81848 576140
rect 81995 576138 81996 576140
rect 82143 576138 82144 576140
rect 82291 576138 82292 576140
rect 82439 576138 82440 576140
rect 82587 576138 82588 576140
rect 82735 576138 82736 576140
rect 82883 576138 82884 576140
rect 83031 576138 83032 576140
rect 83179 576138 83180 576140
rect 83327 576138 83328 576140
rect 83475 576138 83476 576140
rect 83623 576138 83624 576140
rect 83771 576138 83772 576140
rect 83919 576138 83920 576140
rect 84067 576138 84068 576140
rect 84215 576138 84216 576140
rect 84363 576138 84364 576140
rect 84511 576138 84512 576140
rect 84659 576138 84660 576140
rect 84864 576138 84865 576140
rect 85012 576138 85013 576140
rect 85160 576138 85161 576140
rect 85308 576138 85309 576140
rect 85456 576138 85457 576140
rect 85604 576138 85605 576140
rect 85752 576138 85753 576140
rect 85900 576138 85901 576140
rect 86048 576138 86049 576140
rect 86196 576138 86197 576140
rect 86344 576138 86345 576140
rect 86492 576138 86493 576140
rect 86640 576138 86641 576140
rect 86788 576138 86789 576140
rect 86936 576138 86937 576140
rect 87084 576138 87085 576140
rect 87232 576138 87233 576140
rect 87380 576138 87381 576140
rect 87528 576138 87529 576140
rect 87676 576138 87677 576140
rect 87824 576138 87825 576140
rect 87972 576138 87973 576140
rect 88120 576138 88121 576140
rect 88268 576138 88269 576140
rect 88416 576138 88417 576140
rect 88564 576138 88565 576140
rect 88712 576138 88713 576140
rect 88860 576138 88861 576140
rect 89008 576138 89009 576140
rect 89156 576138 89157 576140
rect 89304 576138 89305 576140
rect 89452 576138 89453 576140
rect 89600 576138 89601 576140
rect 89748 576138 89749 576140
rect 89896 576138 89897 576140
rect 90044 576138 90045 576140
rect 90192 576138 90193 576140
rect 80640 576048 80648 576082
rect 80738 576081 80796 576082
rect 80886 576081 80944 576082
rect 81034 576081 81092 576082
rect 81182 576081 81240 576082
rect 81330 576081 81388 576082
rect 81478 576081 81536 576082
rect 81626 576081 81684 576082
rect 81774 576081 81832 576082
rect 81922 576081 81980 576082
rect 82070 576081 82128 576082
rect 82218 576081 82276 576082
rect 82366 576081 82424 576082
rect 82514 576081 82572 576082
rect 82662 576081 82720 576082
rect 82810 576081 82868 576082
rect 82958 576081 83016 576082
rect 83106 576081 83164 576082
rect 83254 576081 83312 576082
rect 83402 576081 83460 576082
rect 83550 576081 83608 576082
rect 83698 576081 83756 576082
rect 83846 576081 83904 576082
rect 83994 576081 84052 576082
rect 84142 576081 84200 576082
rect 84290 576081 84348 576082
rect 84438 576081 84496 576082
rect 84586 576081 84644 576082
rect 84734 576081 84790 576082
rect 84880 576081 84938 576082
rect 85028 576081 85086 576082
rect 85176 576081 85234 576082
rect 85324 576081 85382 576082
rect 85472 576081 85530 576082
rect 85620 576081 85678 576082
rect 85768 576081 85826 576082
rect 85916 576081 85974 576082
rect 86064 576081 86122 576082
rect 86212 576081 86270 576082
rect 86360 576081 86418 576082
rect 86508 576081 86566 576082
rect 86656 576081 86714 576082
rect 86804 576081 86862 576082
rect 86952 576081 87010 576082
rect 87100 576081 87158 576082
rect 87248 576081 87306 576082
rect 87396 576081 87454 576082
rect 87544 576081 87602 576082
rect 87692 576081 87750 576082
rect 87840 576081 87898 576082
rect 87988 576081 88046 576082
rect 88136 576081 88194 576082
rect 88284 576081 88342 576082
rect 88432 576081 88490 576082
rect 88580 576081 88638 576082
rect 88728 576081 88786 576082
rect 88876 576081 88934 576082
rect 89024 576081 89082 576082
rect 89172 576081 89230 576082
rect 89320 576081 89378 576082
rect 89468 576081 89526 576082
rect 89616 576081 89674 576082
rect 89764 576081 89822 576082
rect 89912 576081 89970 576082
rect 90060 576081 90118 576082
rect 90208 576081 90266 576082
rect 80737 576048 80796 576081
rect 80885 576048 80944 576081
rect 81033 576048 81092 576081
rect 81181 576048 81240 576081
rect 81329 576048 81388 576081
rect 81477 576048 81536 576081
rect 81625 576048 81684 576081
rect 81773 576048 81832 576081
rect 81921 576048 81980 576081
rect 82069 576048 82128 576081
rect 82217 576048 82276 576081
rect 82365 576048 82424 576081
rect 82513 576048 82572 576081
rect 82661 576048 82720 576081
rect 82809 576048 82868 576081
rect 82957 576048 83016 576081
rect 83105 576048 83164 576081
rect 83253 576048 83312 576081
rect 83401 576048 83460 576081
rect 83549 576048 83608 576081
rect 83697 576048 83756 576081
rect 83845 576048 83904 576081
rect 83993 576048 84052 576081
rect 84141 576048 84200 576081
rect 84289 576048 84348 576081
rect 84437 576048 84496 576081
rect 84585 576048 84644 576081
rect 80640 576047 80647 576048
rect 82217 576047 82275 576048
rect 82365 576047 82423 576048
rect 82513 576047 82571 576048
rect 82661 576047 82719 576048
rect 82809 576047 82867 576048
rect 82957 576047 83015 576048
rect 83105 576047 83163 576048
rect 83253 576047 83311 576048
rect 83401 576047 83459 576048
rect 83549 576047 83607 576048
rect 83697 576047 83755 576048
rect 83845 576047 83903 576048
rect 83993 576047 84051 576048
rect 84141 576047 84199 576048
rect 84289 576047 84347 576048
rect 84437 576047 84495 576048
rect 84585 576047 84643 576048
rect 84733 576047 84791 576081
rect 84880 576048 84939 576081
rect 85028 576048 85087 576081
rect 85176 576048 85235 576081
rect 85324 576048 85383 576081
rect 85472 576048 85531 576081
rect 85620 576048 85679 576081
rect 85768 576048 85827 576081
rect 85916 576048 85975 576081
rect 86064 576048 86123 576081
rect 86212 576048 86271 576081
rect 86360 576048 86419 576081
rect 86508 576048 86567 576081
rect 86656 576048 86715 576081
rect 86804 576048 86863 576081
rect 86952 576048 87011 576081
rect 87100 576048 87159 576081
rect 87248 576048 87307 576081
rect 87396 576048 87455 576081
rect 87544 576048 87603 576081
rect 87692 576048 87751 576081
rect 87840 576048 87899 576081
rect 87988 576048 88047 576081
rect 88136 576048 88195 576081
rect 88284 576048 88343 576081
rect 88432 576048 88491 576081
rect 88580 576048 88639 576081
rect 88728 576048 88787 576081
rect 88876 576048 88935 576081
rect 89024 576048 89083 576081
rect 89172 576048 89231 576081
rect 89320 576048 89379 576081
rect 89468 576048 89527 576081
rect 89616 576048 89675 576081
rect 89764 576048 89823 576081
rect 89912 576048 89971 576081
rect 90060 576048 90119 576081
rect 90208 576048 90267 576081
rect 84881 576047 84939 576048
rect 85029 576047 85087 576048
rect 88108 575998 88109 576013
rect 88256 575998 88257 576013
rect 88404 575998 88405 576013
rect 88552 575998 88553 576013
rect 88700 575998 88701 576013
rect 88848 575998 88849 576013
rect 88996 575998 88997 576013
rect 89144 575998 89145 576013
rect 80676 575997 80710 575998
rect 80824 575997 80858 575998
rect 80972 575997 81006 575998
rect 81120 575997 81154 575998
rect 81268 575997 81302 575998
rect 81416 575997 81450 575998
rect 81564 575997 81598 575998
rect 81712 575997 81746 575998
rect 81860 575997 81894 575998
rect 82008 575997 82042 575998
rect 82156 575997 82190 575998
rect 82304 575997 82338 575998
rect 82452 575997 82486 575998
rect 82600 575997 82634 575998
rect 82748 575997 82782 575998
rect 82896 575997 82930 575998
rect 83044 575997 83078 575998
rect 83192 575997 83226 575998
rect 83340 575997 83374 575998
rect 83488 575997 83522 575998
rect 83636 575997 83670 575998
rect 83784 575997 83818 575998
rect 83932 575997 83966 575998
rect 84080 575997 84114 575998
rect 84228 575997 84262 575998
rect 84376 575997 84410 575998
rect 84524 575997 84558 575998
rect 84672 575997 84706 575998
rect 80675 575122 80710 575997
rect 80823 575122 80858 575997
rect 80971 575122 81006 575997
rect 81119 575122 81154 575997
rect 81267 575122 81302 575997
rect 81415 575122 81450 575997
rect 81563 575122 81598 575997
rect 81711 575122 81746 575997
rect 81859 575122 81894 575997
rect 82007 575122 82042 575997
rect 82155 575122 82190 575997
rect 82303 575122 82338 575997
rect 82451 575122 82486 575997
rect 82599 575122 82634 575997
rect 82747 575122 82782 575997
rect 82895 575122 82930 575997
rect 83043 575122 83078 575997
rect 83191 575122 83226 575997
rect 83339 575122 83374 575997
rect 83487 575122 83522 575997
rect 83635 575122 83670 575997
rect 83783 575122 83818 575997
rect 83931 575122 83966 575997
rect 84079 575122 84114 575997
rect 84227 575122 84262 575997
rect 84375 575122 84410 575997
rect 84523 575122 84558 575997
rect 84671 575122 84706 575997
rect 84818 575997 84852 575998
rect 84966 575997 85000 575998
rect 85114 575997 85148 575998
rect 85262 575997 85296 575998
rect 85410 575997 85444 575998
rect 85558 575997 85592 575998
rect 85706 575997 85740 575998
rect 85854 575997 85888 575998
rect 86002 575997 86036 575998
rect 86150 575997 86184 575998
rect 86298 575997 86332 575998
rect 86446 575997 86480 575998
rect 86594 575997 86628 575998
rect 86742 575997 86776 575998
rect 86890 575997 86924 575998
rect 87038 575997 87072 575998
rect 87186 575997 87220 575998
rect 87334 575997 87368 575998
rect 87482 575997 87516 575998
rect 87630 575997 87664 575998
rect 87778 575997 87812 575998
rect 87926 575997 87960 575998
rect 88074 575997 88109 575998
rect 88222 575997 88257 575998
rect 88370 575997 88405 575998
rect 88518 575997 88553 575998
rect 88666 575997 88701 575998
rect 88814 575997 88849 575998
rect 88962 575997 88997 575998
rect 89110 575997 89145 575998
rect 89258 575997 89292 575998
rect 89406 575997 89440 575998
rect 89554 575997 89588 575998
rect 89702 575997 89736 575998
rect 89850 575997 89884 575998
rect 89998 575997 90032 575998
rect 84818 575122 84853 575997
rect 84966 575122 85001 575997
rect 85114 575122 85149 575997
rect 85262 575122 85297 575997
rect 85410 575122 85445 575997
rect 85558 575122 85593 575997
rect 85706 575122 85741 575997
rect 85854 575122 85889 575997
rect 86002 575122 86037 575997
rect 86150 575122 86185 575997
rect 86298 575122 86333 575997
rect 86446 575122 86481 575997
rect 86594 575122 86629 575997
rect 86742 575122 86777 575997
rect 86890 575122 86925 575997
rect 87038 575122 87073 575997
rect 87186 575122 87221 575997
rect 87334 575122 87369 575997
rect 87482 575122 87517 575997
rect 87630 575122 87665 575997
rect 87778 575122 87813 575997
rect 87926 575122 87961 575997
rect 88074 575981 88125 575997
rect 88222 575981 88273 575997
rect 88370 575981 88421 575997
rect 88518 575981 88569 575997
rect 88666 575981 88717 575997
rect 88814 575981 88865 575997
rect 88962 575981 89013 575997
rect 89110 575981 89161 575997
rect 88074 575137 88109 575981
rect 88222 575137 88257 575981
rect 88370 575137 88405 575981
rect 88518 575137 88553 575981
rect 88666 575137 88701 575981
rect 88814 575137 88849 575981
rect 88962 575137 88997 575981
rect 89110 575137 89145 575981
rect 88059 575122 88125 575137
rect 88059 575121 88074 575122
rect 88075 575121 88125 575122
rect 88207 575122 88273 575137
rect 88207 575121 88222 575122
rect 88223 575121 88273 575122
rect 88355 575122 88421 575137
rect 88355 575121 88370 575122
rect 88371 575121 88421 575122
rect 88503 575122 88569 575137
rect 88503 575121 88518 575122
rect 88519 575121 88569 575122
rect 88651 575122 88717 575137
rect 88651 575121 88666 575122
rect 88667 575121 88717 575122
rect 88799 575122 88865 575137
rect 88799 575121 88814 575122
rect 88815 575121 88865 575122
rect 88947 575122 89013 575137
rect 88947 575121 88962 575122
rect 88963 575121 89013 575122
rect 89095 575122 89161 575137
rect 89258 575122 89293 575997
rect 89406 575122 89441 575997
rect 89554 575122 89589 575997
rect 89702 575122 89737 575997
rect 89850 575122 89885 575997
rect 89998 575122 90033 575997
rect 136875 575722 136909 576298
rect 136993 575722 137027 576298
rect 137111 575722 137145 576298
rect 137229 575722 137263 576298
rect 137347 575737 137381 576298
rect 137465 575737 137499 576298
rect 137583 575737 137617 576298
rect 137701 575737 137735 576298
rect 137331 575721 137397 575737
rect 137449 575721 137515 575737
rect 137567 575721 137633 575737
rect 137685 575721 137751 575737
rect 137819 575722 137853 576298
rect 137937 575722 137971 576298
rect 138055 575722 138089 576298
rect 138173 575722 138207 576298
rect 138291 575722 138325 576298
rect 138409 575722 138443 576298
rect 138527 575722 138561 576298
rect 138645 575722 138679 576298
rect 138873 575737 138907 576298
rect 138991 575737 139025 576298
rect 139109 575737 139143 576298
rect 139227 575737 139261 576298
rect 139345 575737 139379 576298
rect 139463 575737 139497 576298
rect 139581 575737 139615 576298
rect 139699 575737 139733 576298
rect 139817 575737 139851 576298
rect 139935 575737 139969 576298
rect 140053 575737 140087 576298
rect 140171 575737 140205 576298
rect 140289 575737 140323 576298
rect 140407 575737 140441 576298
rect 140525 575737 140559 576298
rect 140643 575737 140677 576298
rect 143533 576239 143568 577114
rect 143681 576239 143716 577114
rect 143829 576239 143864 577114
rect 143977 576239 144012 577114
rect 144125 576239 144160 577114
rect 144273 576239 144308 577114
rect 144421 576239 144456 577114
rect 144569 576239 144604 577114
rect 144701 577099 144767 577114
rect 144849 577114 144899 577115
rect 144900 577114 144915 577115
rect 144849 577099 144915 577114
rect 144997 577114 145047 577115
rect 145048 577114 145063 577115
rect 144997 577099 145063 577114
rect 145145 577114 145195 577115
rect 145196 577114 145211 577115
rect 145145 577099 145211 577114
rect 145293 577114 145343 577115
rect 145344 577114 145359 577115
rect 145293 577099 145359 577114
rect 145441 577114 145491 577115
rect 145492 577114 145507 577115
rect 145441 577099 145507 577114
rect 145589 577114 145639 577115
rect 145640 577114 145655 577115
rect 145589 577099 145655 577114
rect 145737 577099 145803 577115
rect 144717 576255 144752 577099
rect 144865 576255 144900 577099
rect 145013 576255 145048 577099
rect 145161 576255 145196 577099
rect 145309 576255 145344 577099
rect 145457 576255 145492 577099
rect 145605 576255 145640 577099
rect 145753 576255 145788 577099
rect 144701 576239 144752 576255
rect 144849 576239 144900 576255
rect 144997 576239 145048 576255
rect 145145 576239 145196 576255
rect 145293 576239 145344 576255
rect 145441 576239 145492 576255
rect 145589 576239 145640 576255
rect 145737 576239 145788 576255
rect 143534 576238 143568 576239
rect 143682 576238 143716 576239
rect 143830 576238 143864 576239
rect 143978 576238 144012 576239
rect 144126 576238 144160 576239
rect 144274 576238 144308 576239
rect 144422 576238 144456 576239
rect 144570 576238 144604 576239
rect 144717 576238 144752 576239
rect 144865 576238 144900 576239
rect 145013 576238 145048 576239
rect 145161 576238 145196 576239
rect 145309 576238 145344 576239
rect 145457 576238 145492 576239
rect 145605 576238 145640 576239
rect 145753 576238 145788 576239
rect 144172 576226 144262 576227
rect 144320 576226 144410 576227
rect 144468 576226 144558 576227
rect 144616 576226 144706 576227
rect 144717 576223 144718 576238
rect 144764 576226 144854 576227
rect 144865 576223 144866 576238
rect 144912 576226 145002 576227
rect 145013 576223 145014 576238
rect 145161 576223 145162 576238
rect 145309 576223 145310 576238
rect 145457 576223 145458 576238
rect 145605 576223 145606 576238
rect 145753 576223 145754 576238
rect 145778 576222 145788 576238
rect 145812 576189 145822 577164
rect 146016 577149 146035 577164
rect 146015 577115 146035 577149
rect 146049 577130 146065 577131
rect 146067 577130 146083 577131
rect 146197 577130 146213 577131
rect 146215 577130 146231 577131
rect 146345 577130 146361 577131
rect 146363 577130 146379 577131
rect 146493 577130 146509 577131
rect 146511 577130 146527 577131
rect 146641 577130 146657 577131
rect 146659 577130 146675 577131
rect 146789 577130 146805 577131
rect 146807 577130 146823 577131
rect 146937 577130 146953 577131
rect 146955 577130 146971 577131
rect 147085 577130 147101 577131
rect 147103 577130 147119 577131
rect 147233 577130 147249 577131
rect 147251 577130 147267 577131
rect 147381 577130 147397 577131
rect 147399 577130 147415 577131
rect 147529 577130 147545 577131
rect 147547 577130 147563 577131
rect 147677 577130 147693 577131
rect 147695 577130 147711 577131
rect 147825 577130 147841 577131
rect 147843 577130 147859 577131
rect 147973 577130 147989 577131
rect 147991 577130 148007 577131
rect 148121 577130 148137 577131
rect 148139 577130 148155 577131
rect 148269 577130 148285 577131
rect 148287 577130 148303 577131
rect 148417 577130 148433 577131
rect 148435 577130 148451 577131
rect 146049 577115 146069 577130
rect 146197 577115 146198 577130
rect 146345 577115 146346 577130
rect 146493 577115 146494 577130
rect 146641 577115 146642 577130
rect 146789 577115 146790 577130
rect 146937 577115 146938 577130
rect 147085 577115 147086 577130
rect 147233 577115 147234 577130
rect 147381 577115 147382 577130
rect 147529 577115 147530 577130
rect 147677 577115 147678 577130
rect 147825 577115 147826 577130
rect 147973 577115 147974 577130
rect 148121 577115 148122 577130
rect 148269 577115 148270 577130
rect 148417 577115 148418 577130
rect 145901 577114 145935 577115
rect 146015 577114 146083 577115
rect 146084 577114 146099 577115
rect 145901 576239 145936 577114
rect 145902 576238 145936 576239
rect 146015 577099 146099 577114
rect 146181 577114 146231 577115
rect 146232 577114 146247 577115
rect 146181 577099 146247 577114
rect 146329 577114 146379 577115
rect 146380 577114 146395 577115
rect 146329 577099 146395 577114
rect 146477 577114 146527 577115
rect 146528 577114 146543 577115
rect 146477 577099 146543 577114
rect 146625 577114 146675 577115
rect 146676 577114 146691 577115
rect 146625 577099 146691 577114
rect 146773 577114 146823 577115
rect 146824 577114 146839 577115
rect 146773 577099 146839 577114
rect 146921 577114 146971 577115
rect 146972 577114 146987 577115
rect 146921 577099 146987 577114
rect 147069 577114 147119 577115
rect 147120 577114 147135 577115
rect 147069 577099 147135 577114
rect 147217 577114 147267 577115
rect 147268 577114 147283 577115
rect 147217 577099 147283 577114
rect 147365 577114 147415 577115
rect 147416 577114 147431 577115
rect 147365 577099 147431 577114
rect 147513 577114 147563 577115
rect 147564 577114 147579 577115
rect 147513 577099 147579 577114
rect 147661 577114 147711 577115
rect 147712 577114 147727 577115
rect 147661 577099 147727 577114
rect 147809 577114 147859 577115
rect 147860 577114 147875 577115
rect 147809 577099 147875 577114
rect 147957 577114 148007 577115
rect 148008 577114 148023 577115
rect 147957 577099 148023 577114
rect 148105 577114 148155 577115
rect 148156 577114 148171 577115
rect 148105 577099 148171 577114
rect 148253 577114 148303 577115
rect 148304 577114 148319 577115
rect 148253 577099 148319 577114
rect 148401 577114 148451 577115
rect 148452 577114 148467 577115
rect 148401 577099 148467 577114
rect 148549 577099 148555 577115
rect 146015 576255 146035 577099
rect 146049 576255 146084 577099
rect 146197 576255 146232 577099
rect 146345 576255 146380 577099
rect 146493 576255 146528 577099
rect 146641 576255 146676 577099
rect 146789 576255 146824 577099
rect 146937 576255 146972 577099
rect 147085 576255 147120 577099
rect 147233 576255 147268 577099
rect 147381 576255 147416 577099
rect 147529 576255 147564 577099
rect 147677 576255 147712 577099
rect 147825 576255 147860 577099
rect 147973 576255 148008 577099
rect 148121 576255 148156 577099
rect 148269 576255 148304 577099
rect 148417 576255 148452 577099
rect 146015 576239 146084 576255
rect 146181 576239 146232 576255
rect 146329 576239 146380 576255
rect 146477 576239 146528 576255
rect 146625 576239 146676 576255
rect 146773 576239 146824 576255
rect 146921 576239 146972 576255
rect 147069 576239 147120 576255
rect 147217 576239 147268 576255
rect 147365 576239 147416 576255
rect 147513 576239 147564 576255
rect 147661 576239 147712 576255
rect 147809 576239 147860 576255
rect 147957 576239 148008 576255
rect 148105 576239 148156 576255
rect 148253 576239 148304 576255
rect 148401 576239 148452 576255
rect 148549 576239 148555 576255
rect 146015 576205 146035 576239
rect 146049 576238 146084 576239
rect 146197 576238 146232 576239
rect 146345 576238 146380 576239
rect 146493 576238 146528 576239
rect 146641 576238 146676 576239
rect 146789 576238 146824 576239
rect 146937 576238 146972 576239
rect 147085 576238 147120 576239
rect 147233 576238 147268 576239
rect 147381 576238 147416 576239
rect 147529 576238 147564 576239
rect 147677 576238 147712 576239
rect 147825 576238 147860 576239
rect 147973 576238 148008 576239
rect 148121 576238 148156 576239
rect 148269 576238 148304 576239
rect 148417 576238 148452 576239
rect 146049 576223 146069 576238
rect 146197 576223 146198 576238
rect 146345 576223 146346 576238
rect 146493 576223 146494 576238
rect 146540 576226 146630 576227
rect 146641 576223 146642 576238
rect 146688 576226 146778 576227
rect 146789 576223 146790 576238
rect 146836 576226 146926 576227
rect 146937 576223 146938 576238
rect 146984 576226 147074 576227
rect 147085 576223 147086 576238
rect 147132 576226 147222 576227
rect 147233 576223 147234 576238
rect 147280 576226 147370 576227
rect 147381 576223 147382 576238
rect 147428 576226 147518 576227
rect 147529 576223 147530 576238
rect 147576 576226 147666 576227
rect 147677 576223 147678 576238
rect 147724 576226 147814 576227
rect 147825 576223 147826 576238
rect 147872 576226 147962 576227
rect 147973 576223 147974 576238
rect 148020 576226 148110 576227
rect 148121 576223 148122 576238
rect 148168 576226 148258 576227
rect 148269 576223 148270 576238
rect 148316 576226 148406 576227
rect 148417 576223 148418 576238
rect 148464 576226 148554 576227
rect 146050 576222 146069 576223
rect 146016 576189 146035 576205
rect 144187 576188 144245 576189
rect 144335 576188 144393 576189
rect 144483 576188 144541 576189
rect 144631 576188 144689 576189
rect 144779 576188 144837 576189
rect 144927 576188 144985 576189
rect 146555 576188 146613 576189
rect 146703 576188 146761 576189
rect 146851 576188 146909 576189
rect 146999 576188 147057 576189
rect 147147 576188 147205 576189
rect 147295 576188 147353 576189
rect 147443 576188 147501 576189
rect 147591 576188 147649 576189
rect 147739 576188 147797 576189
rect 147887 576188 147945 576189
rect 148035 576188 148093 576189
rect 148183 576188 148241 576189
rect 148331 576188 148389 576189
rect 148479 576188 148537 576189
rect 143743 576155 143802 576188
rect 143891 576155 143950 576188
rect 144039 576155 144098 576188
rect 144187 576155 144246 576188
rect 144335 576155 144394 576188
rect 144483 576155 144542 576188
rect 144631 576155 144690 576188
rect 144779 576155 144838 576188
rect 144927 576155 144986 576188
rect 145075 576155 145134 576188
rect 145223 576155 145282 576188
rect 145371 576155 145430 576188
rect 145519 576155 145578 576188
rect 145667 576155 145726 576188
rect 145815 576155 145874 576188
rect 145963 576155 146022 576188
rect 146111 576155 146170 576188
rect 146259 576155 146318 576188
rect 146407 576155 146466 576188
rect 146555 576155 146614 576188
rect 146703 576155 146762 576188
rect 146851 576155 146910 576188
rect 146999 576155 147058 576188
rect 147147 576155 147206 576188
rect 147295 576155 147354 576188
rect 147443 576155 147502 576188
rect 147591 576155 147650 576188
rect 147739 576155 147798 576188
rect 147887 576155 147946 576188
rect 148035 576155 148094 576188
rect 148183 576155 148242 576188
rect 148331 576155 148390 576188
rect 148479 576155 148538 576188
rect 143744 576154 143802 576155
rect 143892 576154 143950 576155
rect 144040 576154 144098 576155
rect 144188 576154 144246 576155
rect 144336 576154 144394 576155
rect 144484 576154 144542 576155
rect 144632 576154 144690 576155
rect 144780 576154 144838 576155
rect 144928 576154 144986 576155
rect 145076 576154 145134 576155
rect 145224 576154 145282 576155
rect 145372 576154 145430 576155
rect 145520 576154 145578 576155
rect 145668 576154 145726 576155
rect 145816 576154 145874 576155
rect 145964 576154 146022 576155
rect 146112 576154 146170 576155
rect 146260 576154 146318 576155
rect 146408 576154 146466 576155
rect 146556 576154 146614 576155
rect 146704 576154 146762 576155
rect 146852 576154 146910 576155
rect 147000 576154 147058 576155
rect 147148 576154 147206 576155
rect 147296 576154 147354 576155
rect 147444 576154 147502 576155
rect 147592 576154 147650 576155
rect 147740 576154 147798 576155
rect 147888 576154 147946 576155
rect 148036 576154 148094 576155
rect 148184 576154 148242 576155
rect 148332 576154 148390 576155
rect 148480 576154 148538 576155
rect 143669 576138 143670 576140
rect 143817 576138 143818 576140
rect 143965 576138 143966 576140
rect 144113 576138 144114 576140
rect 144261 576138 144262 576140
rect 144409 576138 144410 576140
rect 144557 576138 144558 576140
rect 144705 576138 144706 576140
rect 144853 576138 144854 576140
rect 145001 576138 145002 576140
rect 145149 576138 145150 576140
rect 145297 576138 145298 576140
rect 145445 576138 145446 576140
rect 145593 576138 145594 576140
rect 145741 576138 145742 576140
rect 145889 576138 145890 576140
rect 146037 576138 146038 576140
rect 146185 576138 146186 576140
rect 146333 576138 146334 576140
rect 146481 576138 146482 576140
rect 146629 576138 146630 576140
rect 146777 576138 146778 576140
rect 146925 576138 146926 576140
rect 147073 576138 147074 576140
rect 147221 576138 147222 576140
rect 147369 576138 147370 576140
rect 147517 576138 147518 576140
rect 147665 576138 147666 576140
rect 147813 576138 147814 576140
rect 147961 576138 147962 576140
rect 148109 576138 148110 576140
rect 148257 576138 148258 576140
rect 148405 576138 148406 576140
rect 148553 576138 148554 576140
rect 143744 576081 143802 576082
rect 143892 576081 143950 576082
rect 144040 576081 144098 576082
rect 144188 576081 144246 576082
rect 144336 576081 144394 576082
rect 144484 576081 144542 576082
rect 144632 576081 144690 576082
rect 144780 576081 144838 576082
rect 144928 576081 144986 576082
rect 145076 576081 145134 576082
rect 145224 576081 145282 576082
rect 145372 576081 145430 576082
rect 145520 576081 145578 576082
rect 145668 576081 145726 576082
rect 145816 576081 145874 576082
rect 145964 576081 146022 576082
rect 146112 576081 146170 576082
rect 146260 576081 146318 576082
rect 146408 576081 146466 576082
rect 146556 576081 146614 576082
rect 146704 576081 146762 576082
rect 146852 576081 146910 576082
rect 147000 576081 147058 576082
rect 147148 576081 147206 576082
rect 147296 576081 147354 576082
rect 147444 576081 147502 576082
rect 147592 576081 147650 576082
rect 147740 576081 147798 576082
rect 147888 576081 147946 576082
rect 148036 576081 148094 576082
rect 148184 576081 148242 576082
rect 148332 576081 148390 576082
rect 148480 576081 148538 576082
rect 143743 576048 143802 576081
rect 143891 576048 143950 576081
rect 144039 576048 144098 576081
rect 144187 576048 144246 576081
rect 144335 576048 144394 576081
rect 144483 576048 144542 576081
rect 144631 576048 144690 576081
rect 144779 576048 144838 576081
rect 144927 576048 144986 576081
rect 145075 576048 145134 576081
rect 145223 576048 145282 576081
rect 145371 576048 145430 576081
rect 145519 576048 145578 576081
rect 145667 576048 145726 576081
rect 145815 576048 145874 576081
rect 145963 576048 146022 576081
rect 146111 576048 146170 576081
rect 146259 576048 146318 576081
rect 146407 576048 146466 576081
rect 146555 576048 146614 576081
rect 146703 576048 146762 576081
rect 146851 576048 146910 576081
rect 146999 576048 147058 576081
rect 147147 576048 147206 576081
rect 147295 576048 147354 576081
rect 147443 576048 147502 576081
rect 147591 576048 147650 576081
rect 147739 576048 147798 576081
rect 147887 576048 147946 576081
rect 148035 576048 148094 576081
rect 148183 576048 148242 576081
rect 148331 576048 148390 576081
rect 148479 576048 148538 576081
rect 144187 576047 144245 576048
rect 144335 576047 144393 576048
rect 144483 576047 144541 576048
rect 144631 576047 144689 576048
rect 144779 576047 144837 576048
rect 144927 576047 144985 576048
rect 146555 576047 146613 576048
rect 146703 576047 146761 576048
rect 146851 576047 146909 576048
rect 146999 576047 147057 576048
rect 147147 576047 147205 576048
rect 147295 576047 147353 576048
rect 147443 576047 147501 576048
rect 147591 576047 147649 576048
rect 147739 576047 147797 576048
rect 147887 576047 147945 576048
rect 148035 576047 148093 576048
rect 148183 576047 148241 576048
rect 148331 576047 148389 576048
rect 148479 576047 148537 576048
rect 145778 575998 145788 576014
rect 143534 575997 143568 575998
rect 143682 575997 143716 575998
rect 143830 575997 143864 575998
rect 143978 575997 144012 575998
rect 144126 575997 144160 575998
rect 144274 575997 144308 575998
rect 144422 575997 144456 575998
rect 144570 575997 144604 575998
rect 144718 575997 144752 575998
rect 144866 575997 144900 575998
rect 145014 575997 145048 575998
rect 145162 575997 145196 575998
rect 145310 575997 145344 575998
rect 145458 575997 145492 575998
rect 145606 575997 145640 575998
rect 145754 575997 145788 575998
rect 138857 575721 138923 575737
rect 138975 575721 139041 575737
rect 139093 575721 139159 575737
rect 139211 575721 139277 575737
rect 139329 575721 139395 575737
rect 139447 575721 139513 575737
rect 139565 575721 139631 575737
rect 139683 575721 139749 575737
rect 139801 575721 139867 575737
rect 139919 575721 139985 575737
rect 140037 575721 140103 575737
rect 140155 575721 140221 575737
rect 140273 575721 140339 575737
rect 140391 575721 140457 575737
rect 140509 575721 140575 575737
rect 140627 575721 140693 575737
rect 137347 575705 137363 575706
rect 137365 575705 137381 575706
rect 137465 575705 137481 575706
rect 137483 575705 137499 575706
rect 137583 575705 137599 575706
rect 137601 575705 137617 575706
rect 137701 575705 137717 575706
rect 137719 575705 137735 575706
rect 138873 575705 138889 575706
rect 138891 575705 138907 575706
rect 138991 575705 139007 575706
rect 139009 575705 139025 575706
rect 139109 575705 139125 575706
rect 139127 575705 139143 575706
rect 139227 575705 139243 575706
rect 139245 575705 139261 575706
rect 139345 575705 139361 575706
rect 139363 575705 139379 575706
rect 139463 575705 139479 575706
rect 139481 575705 139497 575706
rect 139581 575705 139597 575706
rect 139599 575705 139615 575706
rect 139699 575705 139715 575706
rect 139717 575705 139733 575706
rect 139817 575705 139833 575706
rect 139835 575705 139851 575706
rect 139935 575705 139951 575706
rect 139953 575705 139969 575706
rect 140053 575705 140069 575706
rect 140071 575705 140087 575706
rect 140171 575705 140187 575706
rect 140189 575705 140205 575706
rect 140289 575705 140305 575706
rect 140307 575705 140323 575706
rect 140407 575705 140423 575706
rect 140425 575705 140441 575706
rect 140525 575705 140541 575706
rect 140543 575705 140559 575706
rect 140643 575705 140659 575706
rect 140661 575705 140677 575706
rect 143533 575122 143568 575997
rect 143681 575122 143716 575997
rect 143829 575122 143864 575997
rect 143977 575122 144012 575997
rect 144125 575122 144160 575997
rect 144273 575122 144308 575997
rect 144421 575122 144456 575997
rect 144569 575122 144604 575997
rect 144717 575122 144752 575997
rect 144865 575122 144900 575997
rect 145013 575122 145048 575997
rect 145161 575122 145196 575997
rect 145309 575122 145344 575997
rect 145457 575122 145492 575997
rect 145605 575122 145640 575997
rect 145753 575122 145788 575997
rect 89095 575121 89110 575122
rect 89111 575121 89161 575122
rect 88108 575106 88109 575121
rect 88256 575106 88257 575121
rect 88404 575106 88405 575121
rect 88552 575106 88553 575121
rect 88700 575106 88701 575121
rect 88848 575106 88849 575121
rect 88996 575106 88997 575121
rect 89144 575106 89145 575121
rect 145778 575106 145788 575122
rect 88075 575105 88091 575106
rect 88093 575105 88109 575106
rect 88223 575105 88239 575106
rect 88241 575105 88257 575106
rect 88371 575105 88387 575106
rect 88389 575105 88405 575106
rect 88519 575105 88535 575106
rect 88537 575105 88553 575106
rect 88667 575105 88683 575106
rect 88685 575105 88701 575106
rect 88815 575105 88831 575106
rect 88833 575105 88849 575106
rect 88963 575105 88979 575106
rect 88981 575105 88997 575106
rect 89111 575105 89127 575106
rect 89129 575105 89145 575106
rect 145812 575072 145822 576047
rect 146016 576031 146035 576047
rect 145902 575997 145936 575998
rect 145901 575122 145936 575997
rect 146015 575087 146035 576031
rect 146050 575998 146069 576014
rect 146050 575997 146084 575998
rect 146198 575997 146232 575998
rect 146346 575997 146380 575998
rect 146494 575997 146528 575998
rect 146642 575997 146676 575998
rect 146790 575997 146824 575998
rect 146938 575997 146972 575998
rect 147086 575997 147120 575998
rect 147234 575997 147268 575998
rect 147382 575997 147416 575998
rect 147530 575997 147564 575998
rect 147678 575997 147712 575998
rect 147826 575997 147860 575998
rect 147974 575997 148008 575998
rect 148122 575997 148156 575998
rect 148270 575997 148304 575998
rect 148418 575997 148452 575998
rect 146049 575122 146084 575997
rect 146197 575122 146232 575997
rect 146345 575122 146380 575997
rect 146493 575122 146528 575997
rect 146641 575122 146676 575997
rect 146789 575122 146824 575997
rect 146937 575122 146972 575997
rect 147085 575122 147120 575997
rect 147233 575122 147268 575997
rect 147381 575122 147416 575997
rect 147529 575122 147564 575997
rect 147677 575122 147712 575997
rect 147825 575122 147860 575997
rect 147973 575122 148008 575997
rect 148121 575122 148156 575997
rect 148269 575122 148304 575997
rect 148417 575122 148452 575997
rect 146049 575121 146069 575122
rect 146050 575106 146069 575121
rect 146016 575072 146035 575087
rect 128306 556573 128322 557250
rect 128294 556545 128322 556573
rect 128294 556517 128334 556545
rect 128306 556489 128334 556517
rect 164480 549157 164486 549162
rect 164474 549150 164479 549156
rect 164474 547596 164479 547602
rect 164480 547590 164486 547595
<< poly >>
rect 129936 568408 129996 568424
rect 129936 568374 129952 568408
rect 129986 568406 129996 568408
rect 130638 568410 130698 568426
rect 130638 568406 130648 568410
rect 129986 568376 130648 568406
rect 130682 568376 130698 568410
rect 129986 568374 129996 568376
rect 129936 568358 129996 568374
rect 130638 568360 130698 568376
rect 129906 556348 129966 556364
rect 129906 556314 129922 556348
rect 129956 556346 129966 556348
rect 130608 556346 130668 556362
rect 129956 556316 130618 556346
rect 129956 556314 129966 556316
rect 129906 556298 129966 556314
rect 130608 556312 130618 556316
rect 130652 556312 130668 556346
rect 130608 556296 130668 556312
rect 130042 483716 130102 483732
rect 130042 483682 130058 483716
rect 130092 483714 130102 483716
rect 130744 483718 130804 483734
rect 130744 483714 130754 483718
rect 130092 483684 130754 483714
rect 130788 483684 130804 483718
rect 130092 483682 130102 483684
rect 130042 483666 130102 483682
rect 130744 483668 130804 483684
<< polycont >>
rect 129952 568374 129986 568408
rect 130648 568376 130682 568410
rect 129922 556314 129956 556348
rect 130618 556312 130652 556346
rect 130058 483682 130092 483716
rect 130754 483684 130788 483718
<< locali >>
rect 121460 580842 123290 580848
rect 121460 580674 129849 580842
rect 121460 579148 121662 580674
rect 123066 579148 129849 580674
rect 121460 578952 129849 579148
rect 121460 576732 123290 576738
rect 121460 576564 129625 576732
rect 121460 575038 121662 576564
rect 123066 575038 129625 576564
rect 121460 574842 129625 575038
rect 121460 572800 123290 572806
rect 121460 572632 129687 572800
rect 121460 571106 121662 572632
rect 123066 571106 129687 572632
rect 121460 570910 129687 571106
rect 121460 568958 123290 568964
rect 121460 568790 129687 568958
rect 121460 567264 121662 568790
rect 123066 568594 129687 568790
rect 123066 568408 129986 568594
rect 130865 568569 131088 572491
rect 145812 569815 146035 583940
rect 186090 580658 187920 580664
rect 186090 580490 194236 580658
rect 186090 578964 186292 580490
rect 187696 578964 194236 580490
rect 186090 578768 194236 578964
rect 186060 576898 187890 576904
rect 186060 576730 194206 576898
rect 186060 575204 186262 576730
rect 187666 575204 194206 576730
rect 186060 575008 194206 575204
rect 186060 573258 187890 573264
rect 186060 573090 194206 573258
rect 186060 571564 186262 573090
rect 187666 571564 194206 573090
rect 186060 571368 194206 571564
rect 130649 568568 131088 568569
rect 123066 568374 129952 568408
rect 123066 568186 129986 568374
rect 130648 568410 131088 568568
rect 130682 568376 131088 568410
rect 130648 568344 131088 568376
rect 130649 568343 131088 568344
rect 123066 567264 129687 568186
rect 121460 567068 129687 567264
rect 121446 557010 123276 557016
rect 121446 556842 129687 557010
rect 121446 555316 121648 556842
rect 123052 556536 129687 556842
rect 123052 556348 129956 556536
rect 130619 556378 131058 556379
rect 123052 556314 129922 556348
rect 123052 556128 129956 556314
rect 130618 556346 131058 556378
rect 130652 556312 131058 556346
rect 130618 556154 131058 556312
rect 130619 556153 131058 556154
rect 123052 555316 129687 556128
rect 121446 555120 129687 555316
rect 121460 553466 123290 553472
rect 121460 553298 129701 553466
rect 121460 551772 121662 553298
rect 123066 551772 129701 553298
rect 130835 552629 131058 556153
rect 186060 553450 187890 553456
rect 186060 553282 194206 553450
rect 121460 551576 129701 551772
rect 186060 551756 186262 553282
rect 187666 551756 194206 553282
rect 186060 551560 194206 551756
rect 121460 549862 123290 549868
rect 121460 549694 129701 549862
rect 121460 548168 121662 549694
rect 123066 548168 129701 549694
rect 121460 547972 129701 548168
rect 186060 549406 187890 549412
rect 186060 549238 194206 549406
rect 186060 547712 186262 549238
rect 187666 547712 194206 549238
rect 186060 547516 194206 547712
rect 121460 545930 123290 545936
rect 121460 545762 129715 545930
rect 121460 544236 121662 545762
rect 123066 544236 129715 545762
rect 121460 544040 129715 544236
rect 186060 545768 187890 545774
rect 186060 545600 194206 545768
rect 186060 544074 186262 545600
rect 187666 544074 194206 545600
rect 186060 543878 194206 544074
rect 121460 495466 123290 495472
rect 121460 495298 130037 495466
rect 121460 493772 121662 495298
rect 123066 493772 130037 495298
rect 121460 493576 130037 493772
rect 121460 491534 123290 491540
rect 121460 491366 129980 491534
rect 121460 489840 121662 491366
rect 123066 489840 129980 491366
rect 121460 489650 129980 489840
rect 121460 489644 123866 489650
rect 121460 487930 123290 487936
rect 121460 487762 129983 487930
rect 121460 486236 121662 487762
rect 123066 486236 129983 487762
rect 121460 486040 129983 486236
rect 121432 484342 123262 484348
rect 121432 484174 129955 484342
rect 121432 482648 121634 484174
rect 123038 483902 129955 484174
rect 123038 483716 130092 483902
rect 130971 483877 131194 487315
rect 130755 483876 131194 483877
rect 123038 483682 130058 483716
rect 123038 483494 130092 483682
rect 130754 483718 131194 483876
rect 130788 483684 131194 483718
rect 130754 483652 131194 483684
rect 130755 483651 131194 483652
rect 123038 482648 129955 483494
rect 121432 482452 129955 482648
<< viali >>
rect 121662 579148 123066 580674
rect 121662 575038 123066 576564
rect 121662 571106 123066 572632
rect 121662 567264 123066 568790
rect 186292 578964 187696 580490
rect 186262 575204 187666 576730
rect 186262 571564 187666 573090
rect 121648 555316 123052 556842
rect 121662 551772 123066 553298
rect 186262 551756 187666 553282
rect 121662 548168 123066 549694
rect 186262 547712 187666 549238
rect 121662 544236 123066 545762
rect 186262 544074 187666 545600
rect 121662 493772 123066 495298
rect 121662 489840 123066 491366
rect 121662 486236 123066 487762
rect 121634 482648 123038 484174
<< metal1 >>
rect 121598 580674 123138 580726
rect 121598 580668 121662 580674
rect 123066 580668 123138 580674
rect 121598 579132 121648 580668
rect 123096 579132 123138 580668
rect 121598 579082 123138 579132
rect 186228 580490 187768 580542
rect 186228 580484 186292 580490
rect 187696 580484 187768 580490
rect 186228 578948 186278 580484
rect 187726 578948 187768 580484
rect 186228 578898 187768 578948
rect 186198 576730 187738 576782
rect 186198 576724 186262 576730
rect 187666 576724 187738 576730
rect 121598 576564 123138 576616
rect 121598 576558 121662 576564
rect 123066 576558 123138 576564
rect 121598 575022 121648 576558
rect 123096 575022 123138 576558
rect 186198 575188 186248 576724
rect 187696 575188 187738 576724
rect 186198 575138 187738 575188
rect 121598 574972 123138 575022
rect 186198 573090 187738 573142
rect 186198 573084 186262 573090
rect 187666 573084 187738 573090
rect 121598 572632 123138 572684
rect 121598 572626 121662 572632
rect 123066 572626 123138 572632
rect 121598 571090 121648 572626
rect 123096 571090 123138 572626
rect 186198 571548 186248 573084
rect 187696 571548 187738 573084
rect 186198 571498 187738 571548
rect 121598 571040 123138 571090
rect 121598 568790 123138 568842
rect 121598 568784 121662 568790
rect 123066 568784 123138 568790
rect 121598 567248 121648 568784
rect 123096 567248 123138 568784
rect 121598 567198 123138 567248
rect 121584 556842 123124 556894
rect 121584 556836 121648 556842
rect 123052 556836 123124 556842
rect 121584 555300 121634 556836
rect 123082 555300 123124 556836
rect 121584 555250 123124 555300
rect 121598 553298 123138 553350
rect 121598 553292 121662 553298
rect 123066 553292 123138 553298
rect 121598 551756 121648 553292
rect 123096 551756 123138 553292
rect 121598 551706 123138 551756
rect 186198 553282 187738 553334
rect 186198 553276 186262 553282
rect 187666 553276 187738 553282
rect 186198 551740 186248 553276
rect 187696 551740 187738 553276
rect 186198 551690 187738 551740
rect 121598 549694 123138 549746
rect 121598 549688 121662 549694
rect 123066 549688 123138 549694
rect 121598 548152 121648 549688
rect 123096 548152 123138 549688
rect 121598 548102 123138 548152
rect 186198 549238 187738 549290
rect 186198 549232 186262 549238
rect 187666 549232 187738 549238
rect 186198 547696 186248 549232
rect 187696 547696 187738 549232
rect 186198 547646 187738 547696
rect 121598 545762 123138 545814
rect 121598 545756 121662 545762
rect 123066 545756 123138 545762
rect 121598 544220 121648 545756
rect 123096 544220 123138 545756
rect 121598 544170 123138 544220
rect 186198 545600 187738 545652
rect 186198 545594 186262 545600
rect 187666 545594 187738 545600
rect 186198 544058 186248 545594
rect 187696 544058 187738 545594
rect 186198 544008 187738 544058
rect 121598 495298 123138 495350
rect 121598 495292 121662 495298
rect 123066 495292 123138 495298
rect 121598 493756 121648 495292
rect 123096 493756 123138 495292
rect 121598 493706 123138 493756
rect 121598 491366 123138 491418
rect 121598 491360 121662 491366
rect 123066 491360 123138 491366
rect 121598 489824 121648 491360
rect 123096 489824 123138 491360
rect 121598 489774 123138 489824
rect 121598 487762 123138 487814
rect 121598 487756 121662 487762
rect 123066 487756 123138 487762
rect 121598 486220 121648 487756
rect 123096 486220 123138 487756
rect 121598 486170 123138 486220
rect 121570 484174 123110 484226
rect 121570 484168 121634 484174
rect 123038 484168 123110 484174
rect 121570 482632 121620 484168
rect 123068 482632 123110 484168
rect 121570 482582 123110 482632
<< via1 >>
rect 121648 579148 121662 580668
rect 121662 579148 123066 580668
rect 123066 579148 123096 580668
rect 121648 579132 123096 579148
rect 186278 578964 186292 580484
rect 186292 578964 187696 580484
rect 187696 578964 187726 580484
rect 186278 578948 187726 578964
rect 121648 575038 121662 576558
rect 121662 575038 123066 576558
rect 123066 575038 123096 576558
rect 121648 575022 123096 575038
rect 186248 575204 186262 576724
rect 186262 575204 187666 576724
rect 187666 575204 187696 576724
rect 186248 575188 187696 575204
rect 121648 571106 121662 572626
rect 121662 571106 123066 572626
rect 123066 571106 123096 572626
rect 121648 571090 123096 571106
rect 186248 571564 186262 573084
rect 186262 571564 187666 573084
rect 187666 571564 187696 573084
rect 186248 571548 187696 571564
rect 121648 567264 121662 568784
rect 121662 567264 123066 568784
rect 123066 567264 123096 568784
rect 121648 567248 123096 567264
rect 121634 555316 121648 556836
rect 121648 555316 123052 556836
rect 123052 555316 123082 556836
rect 121634 555300 123082 555316
rect 121648 551772 121662 553292
rect 121662 551772 123066 553292
rect 123066 551772 123096 553292
rect 121648 551756 123096 551772
rect 186248 551756 186262 553276
rect 186262 551756 187666 553276
rect 187666 551756 187696 553276
rect 186248 551740 187696 551756
rect 121648 548168 121662 549688
rect 121662 548168 123066 549688
rect 123066 548168 123096 549688
rect 121648 548152 123096 548168
rect 186248 547712 186262 549232
rect 186262 547712 187666 549232
rect 187666 547712 187696 549232
rect 186248 547696 187696 547712
rect 121648 544236 121662 545756
rect 121662 544236 123066 545756
rect 123066 544236 123096 545756
rect 121648 544220 123096 544236
rect 186248 544074 186262 545594
rect 186262 544074 187666 545594
rect 187666 544074 187696 545594
rect 186248 544058 187696 544074
rect 121648 493772 121662 495292
rect 121662 493772 123066 495292
rect 123066 493772 123096 495292
rect 121648 493756 123096 493772
rect 121648 489840 121662 491360
rect 121662 489840 123066 491360
rect 123066 489840 123096 491360
rect 121648 489824 123096 489840
rect 121648 486236 121662 487756
rect 121662 486236 123066 487756
rect 123066 486236 123096 487756
rect 121648 486220 123096 486236
rect 121620 482648 121634 484168
rect 121634 482648 123038 484168
rect 123038 482648 123068 484168
rect 121620 482632 123068 482648
<< metal2 >>
rect 51490 640921 58420 640930
rect 51490 597173 58420 633991
rect 66834 597173 67014 597178
rect 195514 597173 195680 597180
rect 51490 597000 195680 597173
rect 51490 596188 195687 597000
rect 51490 529437 58420 596188
rect 66834 592876 67014 596188
rect 131176 593004 131349 596188
rect 195514 591943 195687 596188
rect 121518 580710 123212 580798
rect 121518 579090 121604 580710
rect 123124 579090 123212 580710
rect 121518 579002 123212 579090
rect 186148 580526 187842 580614
rect 186148 578906 186234 580526
rect 187754 578906 187842 580526
rect 186148 578818 187842 578906
rect 186118 576766 187812 576854
rect 121518 576600 123212 576688
rect 121518 574980 121604 576600
rect 123124 574980 123212 576600
rect 186118 575146 186204 576766
rect 187724 575146 187812 576766
rect 186118 575058 187812 575146
rect 121518 574892 123212 574980
rect 186118 573126 187812 573214
rect 121518 572668 123212 572756
rect 121518 571048 121604 572668
rect 123124 571048 123212 572668
rect 186118 571506 186204 573126
rect 187724 571506 187812 573126
rect 186118 571418 187812 571506
rect 121518 570960 123212 571048
rect 121518 568826 123212 568914
rect 121518 567206 121604 568826
rect 123124 567206 123212 568826
rect 121518 567118 123212 567206
rect 121504 556878 123198 556966
rect 121504 555258 121590 556878
rect 123110 555258 123198 556878
rect 128294 556517 128306 557250
rect 121504 555170 123198 555258
rect 121518 553334 123212 553422
rect 121518 551714 121604 553334
rect 123124 551714 123212 553334
rect 121518 551626 123212 551714
rect 186118 553318 187812 553406
rect 186118 551698 186204 553318
rect 187724 551698 187812 553318
rect 186118 551610 187812 551698
rect 121518 549730 123212 549818
rect 121518 548110 121604 549730
rect 123124 548110 123212 549730
rect 121518 548022 123212 548110
rect 186118 549274 187812 549362
rect 186118 547654 186204 549274
rect 187724 547654 187812 549274
rect 186118 547566 187812 547654
rect 121518 545798 123212 545886
rect 121518 544178 121604 545798
rect 123124 544178 123212 545798
rect 121518 544090 123212 544178
rect 186118 545636 187812 545724
rect 186118 544016 186204 545636
rect 187724 544016 187812 545636
rect 186118 543928 187812 544016
rect 66822 529437 66995 532135
rect 131160 529437 131333 533807
rect 195498 529437 195671 532271
rect 51490 528452 195671 529437
rect 51490 511471 58420 528452
rect 195498 528448 195671 528452
rect 51490 510486 131530 511471
rect 51490 443429 58420 510486
rect 66682 507929 66855 510486
rect 131310 507468 131483 510486
rect 121518 495334 123212 495422
rect 121518 493714 121604 495334
rect 123124 493714 123212 495334
rect 121518 493626 123212 493714
rect 121518 491402 123212 491490
rect 121518 489782 121604 491402
rect 123124 489782 123212 491402
rect 121518 489694 123212 489782
rect 121518 487798 123212 487886
rect 121518 486178 121604 487798
rect 123124 486178 123212 487798
rect 121518 486090 123212 486178
rect 121490 484210 123184 484298
rect 121490 482590 121576 484210
rect 123096 482590 123184 484210
rect 121490 482502 123184 482590
rect 66666 443429 66839 447381
rect 51490 442450 66839 443429
rect 51490 442444 66708 442450
rect 51490 442436 58420 442444
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 51490 633991 58420 640921
rect 121604 580668 123124 580710
rect 121604 579132 121648 580668
rect 121648 579132 123096 580668
rect 123096 579132 123124 580668
rect 121604 579090 123124 579132
rect 186234 580484 187754 580526
rect 186234 578948 186278 580484
rect 186278 578948 187726 580484
rect 187726 578948 187754 580484
rect 186234 578906 187754 578948
rect 121604 576558 123124 576600
rect 121604 575022 121648 576558
rect 121648 575022 123096 576558
rect 123096 575022 123124 576558
rect 121604 574980 123124 575022
rect 186204 576724 187724 576766
rect 186204 575188 186248 576724
rect 186248 575188 187696 576724
rect 187696 575188 187724 576724
rect 186204 575146 187724 575188
rect 121604 572626 123124 572668
rect 121604 571090 121648 572626
rect 121648 571090 123096 572626
rect 123096 571090 123124 572626
rect 121604 571048 123124 571090
rect 186204 573084 187724 573126
rect 186204 571548 186248 573084
rect 186248 571548 187696 573084
rect 187696 571548 187724 573084
rect 186204 571506 187724 571548
rect 121604 568784 123124 568826
rect 121604 567248 121648 568784
rect 121648 567248 123096 568784
rect 123096 567248 123124 568784
rect 121604 567206 123124 567248
rect 121590 556836 123110 556878
rect 121590 555300 121634 556836
rect 121634 555300 123082 556836
rect 123082 555300 123110 556836
rect 121590 555258 123110 555300
rect 121604 553292 123124 553334
rect 121604 551756 121648 553292
rect 121648 551756 123096 553292
rect 123096 551756 123124 553292
rect 121604 551714 123124 551756
rect 186204 553276 187724 553318
rect 186204 551740 186248 553276
rect 186248 551740 187696 553276
rect 187696 551740 187724 553276
rect 186204 551698 187724 551740
rect 121604 549688 123124 549730
rect 121604 548152 121648 549688
rect 121648 548152 123096 549688
rect 123096 548152 123124 549688
rect 121604 548110 123124 548152
rect 186204 549232 187724 549274
rect 186204 547696 186248 549232
rect 186248 547696 187696 549232
rect 187696 547696 187724 549232
rect 186204 547654 187724 547696
rect 121604 545756 123124 545798
rect 121604 544220 121648 545756
rect 121648 544220 123096 545756
rect 123096 544220 123124 545756
rect 121604 544178 123124 544220
rect 186204 545594 187724 545636
rect 186204 544058 186248 545594
rect 186248 544058 187696 545594
rect 187696 544058 187724 545594
rect 186204 544016 187724 544058
rect 121604 495292 123124 495334
rect 121604 493756 121648 495292
rect 121648 493756 123096 495292
rect 123096 493756 123124 495292
rect 121604 493714 123124 493756
rect 121604 491360 123124 491402
rect 121604 489824 121648 491360
rect 121648 489824 123096 491360
rect 123096 489824 123124 491360
rect 121604 489782 123124 489824
rect 121604 487756 123124 487798
rect 121604 486220 121648 487756
rect 121648 486220 123096 487756
rect 123096 486220 123124 487756
rect 121604 486178 123124 486220
rect 121576 484168 123096 484210
rect 121576 482632 121620 484168
rect 121620 482632 123068 484168
rect 123068 482632 123096 484168
rect 121576 482590 123096 482632
<< metal3 >>
rect 16194 702300 21194 704800
rect -800 680242 1700 685242
rect 68194 663497 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 671294 515394 704800
rect 520594 669112 525394 704800
rect 566594 698484 571594 704800
rect 566594 693478 571594 693484
rect 582300 682980 584800 682984
rect 563698 677984 565634 682980
rect 570630 677984 584800 682980
rect 51490 656567 73409 663497
rect -800 643842 1660 648642
rect 51490 640926 58420 656567
rect 51485 640921 58425 640926
rect -800 633842 1660 638642
rect 51485 633991 51490 640921
rect 58420 633991 58425 640921
rect 582340 639784 584800 644584
rect 51485 633986 58425 633991
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 114778 581446 117484 581712
rect 114778 579580 115042 581446
rect 114748 579372 115042 579580
rect 117144 579372 117484 581446
rect 114748 579122 117484 579372
rect 121402 580826 123328 580928
rect 40405 565352 42711 565357
rect 34738 565351 42712 565352
rect 34738 564242 40405 565351
rect -800 563045 40405 564242
rect 42711 563045 42712 565351
rect 114748 563203 117454 579122
rect 121402 578974 121488 580826
rect 123240 578974 123328 580826
rect 186032 580642 187958 580744
rect 121402 578872 123328 578974
rect 181481 580321 183043 580322
rect 181481 578761 181482 580321
rect 183042 578761 183043 580321
rect 121402 576716 123328 576818
rect 121402 574864 121488 576716
rect 123240 574864 123328 576716
rect 121402 574762 123328 574864
rect 121402 572784 123328 572886
rect 121402 570932 121488 572784
rect 123240 570932 123328 572784
rect 121402 570830 123328 570932
rect 121402 568942 123328 569044
rect 121402 567090 121488 568942
rect 123240 567090 123328 568942
rect 121402 566988 123328 567090
rect -800 563044 42712 563045
rect -800 563039 42711 563044
rect -800 561975 42616 563039
rect -800 559669 40139 561975
rect 42445 559669 42616 561975
rect 114742 560497 114748 563203
rect 117454 560497 117460 563203
rect -800 559442 42616 559669
rect 34738 559388 37046 559442
rect 114748 557651 117454 560497
rect 114748 556994 123439 557651
rect 114748 555142 121474 556994
rect 123226 555142 123439 556994
rect 114748 554945 123439 555142
rect -800 549442 36578 554242
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 28448 480757 36578 549442
rect 101096 553626 123580 553858
rect 101096 551460 101430 553626
rect 103522 553450 123580 553626
rect 103522 551598 121488 553450
rect 123240 551598 123580 553450
rect 181481 553401 183043 578761
rect 186032 578790 186118 580642
rect 187870 578790 187958 580642
rect 186032 578688 187958 578790
rect 186002 576882 187928 576984
rect 186002 575030 186088 576882
rect 187840 575030 187928 576882
rect 186002 574928 187928 575030
rect 186002 573242 187928 573344
rect 186002 571390 186088 573242
rect 187840 571390 187928 573242
rect 186002 571288 187928 571390
rect 186002 553434 187928 553536
rect 186002 553401 186088 553434
rect 181481 551839 186088 553401
rect 187840 553401 187928 553434
rect 103522 551460 123580 551598
rect 186002 551582 186088 551839
rect 187840 551839 188155 553401
rect 187840 551582 187928 551839
rect 186002 551480 187928 551582
rect 101096 551242 123580 551460
rect 101096 535208 103712 551242
rect 487747 550562 487753 566680
rect 503871 555362 559864 566680
rect 503871 550562 584800 555362
rect 121402 549846 123328 549948
rect 106354 549784 109178 549804
rect 121402 549784 121488 549846
rect 106354 549502 121488 549784
rect 123240 549784 123328 549846
rect 106354 547336 106858 549502
rect 108950 547994 121488 549502
rect 123240 547994 123651 549784
rect 186002 549390 187928 549492
rect 186002 549157 186088 549390
rect 108950 547336 123651 547994
rect 164479 549156 186088 549157
rect 164479 547596 164480 549156
rect 166040 547596 186088 549156
rect 164479 547595 186088 547596
rect 186002 547538 186088 547595
rect 187840 547538 187928 549390
rect 186002 547436 187928 547538
rect 106354 547098 123651 547336
rect 121110 545914 123476 546188
rect 121110 545514 121488 545914
rect 111782 545174 121488 545514
rect 111782 542488 112142 545174
rect 114828 544062 121488 545174
rect 123240 545514 123476 545914
rect 186002 545752 187928 545854
rect 123240 544062 123493 545514
rect 114828 542488 123493 544062
rect 186002 543900 186088 545752
rect 187840 543900 187928 545752
rect 186002 543798 187928 543900
rect 111782 541920 123493 542488
rect 527394 540562 584800 545362
rect 101096 532592 114074 535208
rect 111458 496176 114074 532592
rect 103002 494539 104586 494540
rect 102997 492957 103003 494539
rect 104585 492957 104591 494539
rect 111458 493560 117808 496176
rect 103002 487634 104586 492957
rect 115192 492020 117808 493560
rect 121402 495450 123328 495552
rect 121402 493598 121488 495450
rect 123240 493598 123328 495450
rect 121402 493496 123328 493598
rect 115192 491620 123290 492020
rect 115192 491518 123328 491620
rect 115192 489666 121488 491518
rect 123240 489666 123328 491518
rect 115192 489564 123328 489666
rect 115192 489404 123290 489564
rect 121402 487914 123328 488016
rect 121402 487634 121488 487914
rect 103002 486062 121488 487634
rect 123240 486062 123328 487914
rect 103002 486050 123328 486062
rect 121402 485960 123328 486050
rect 121374 484326 123300 484428
rect 121374 482474 121460 484326
rect 123212 482474 123300 484326
rect 121374 482372 123300 482474
rect 28448 478451 33509 480757
rect 35815 478451 36578 480757
rect 28448 477029 36578 478451
rect 28448 474723 29695 477029
rect 32001 474723 36578 477029
rect 28448 474506 36578 474723
rect 527394 481837 543844 540562
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect 527394 463931 543844 465387
rect 539044 463930 543844 463931
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 522540 235230 584800 240030
rect 520920 225230 584800 230030
rect -800 214888 40066 219688
rect -800 204888 47926 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 538388 146830 584800 151630
rect 533702 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 566594 693484 571594 698484
rect 565634 677984 570630 682980
rect 115042 579372 117144 581446
rect 40405 563045 42711 565351
rect 121488 580710 123240 580826
rect 121488 579090 121604 580710
rect 121604 579090 123124 580710
rect 123124 579090 123240 580710
rect 121488 578974 123240 579090
rect 181482 578761 183042 580321
rect 121488 576600 123240 576716
rect 121488 574980 121604 576600
rect 121604 574980 123124 576600
rect 123124 574980 123240 576600
rect 121488 574864 123240 574980
rect 121488 572668 123240 572784
rect 121488 571048 121604 572668
rect 121604 571048 123124 572668
rect 123124 571048 123240 572668
rect 121488 570932 123240 571048
rect 121488 568826 123240 568942
rect 121488 567206 121604 568826
rect 121604 567206 123124 568826
rect 123124 567206 123240 568826
rect 121488 567090 123240 567206
rect 40139 559669 42445 561975
rect 114748 560497 117454 563203
rect 121474 556878 123226 556994
rect 121474 555258 121590 556878
rect 121590 555258 123110 556878
rect 123110 555258 123226 556878
rect 121474 555142 123226 555258
rect 101430 551460 103522 553626
rect 121488 553334 123240 553450
rect 121488 551714 121604 553334
rect 121604 551714 123124 553334
rect 123124 551714 123240 553334
rect 121488 551598 123240 551714
rect 186118 580526 187870 580642
rect 186118 578906 186234 580526
rect 186234 578906 187754 580526
rect 187754 578906 187870 580526
rect 186118 578790 187870 578906
rect 186088 576766 187840 576882
rect 186088 575146 186204 576766
rect 186204 575146 187724 576766
rect 187724 575146 187840 576766
rect 186088 575030 187840 575146
rect 186088 573126 187840 573242
rect 186088 571506 186204 573126
rect 186204 571506 187724 573126
rect 187724 571506 187840 573126
rect 186088 571390 187840 571506
rect 186088 553318 187840 553434
rect 186088 551698 186204 553318
rect 186204 551698 187724 553318
rect 187724 551698 187840 553318
rect 186088 551582 187840 551698
rect 487753 550562 503871 566680
rect 121488 549730 123240 549846
rect 106858 547336 108950 549502
rect 121488 548110 121604 549730
rect 121604 548110 123124 549730
rect 123124 548110 123240 549730
rect 121488 547994 123240 548110
rect 186088 549274 187840 549390
rect 164480 547596 166040 549156
rect 186088 547654 186204 549274
rect 186204 547654 187724 549274
rect 187724 547654 187840 549274
rect 186088 547538 187840 547654
rect 121488 545798 123240 545914
rect 112142 542488 114828 545174
rect 121488 544178 121604 545798
rect 121604 544178 123124 545798
rect 123124 544178 123240 545798
rect 121488 544062 123240 544178
rect 186088 545636 187840 545752
rect 186088 544016 186204 545636
rect 186204 544016 187724 545636
rect 187724 544016 187840 545636
rect 186088 543900 187840 544016
rect 103003 492957 104585 494539
rect 121488 495334 123240 495450
rect 121488 493714 121604 495334
rect 121604 493714 123124 495334
rect 123124 493714 123240 495334
rect 121488 493598 123240 493714
rect 121488 491402 123240 491518
rect 121488 489782 121604 491402
rect 121604 489782 123124 491402
rect 123124 489782 123240 491402
rect 121488 489666 123240 489782
rect 121488 487798 123240 487914
rect 121488 486178 121604 487798
rect 121604 486178 123124 487798
rect 123124 486178 123240 487798
rect 121488 486062 123240 486178
rect 121460 484210 123212 484326
rect 121460 482590 121576 484210
rect 121576 482590 123096 484210
rect 123096 482590 123212 484210
rect 121460 482474 123212 482590
rect 33509 478451 35815 480757
rect 29695 474723 32001 477029
rect 527394 465387 543844 481837
<< metal4 >>
rect 565842 698484 573002 699242
rect 565842 696801 566594 698484
rect 533961 696547 566594 696801
rect 532969 693484 566594 696547
rect 571594 693484 573002 698484
rect 532969 692952 573002 693484
rect 532969 692919 572777 692952
rect 381275 649115 385157 649319
rect 532969 649115 543927 692919
rect 381275 648805 543927 649115
rect 377935 638157 543927 648805
rect 563013 682980 573679 683257
rect 563013 677984 565634 682980
rect 570630 677984 573679 682980
rect 377935 583350 388409 638157
rect 563013 593207 573679 677984
rect 114748 581446 117572 581800
rect 114748 580600 115042 581446
rect 93232 579372 115042 580600
rect 117144 580600 117572 581446
rect 121198 580826 123530 581072
rect 121198 580600 121488 580826
rect 117144 579372 121488 580600
rect 93232 579016 121488 579372
rect 121198 578974 121488 579016
rect 123240 578974 123530 580826
rect 185828 580642 188160 580888
rect 181352 580322 183222 580516
rect 185828 580416 186118 580642
rect 185814 580322 186118 580416
rect 121198 578694 123530 578974
rect 157570 580321 186118 580322
rect 157570 578761 181482 580321
rect 183042 578790 186118 580321
rect 187870 580322 188160 580642
rect 187870 578790 188755 580322
rect 221908 579468 388409 583350
rect 448623 592989 452505 593117
rect 454221 592989 573679 593207
rect 448623 591427 573679 592989
rect 448623 584769 573807 591427
rect 183042 578761 188755 578790
rect 157570 578760 188755 578761
rect 185828 578510 188160 578760
rect 121198 576716 123530 576962
rect 121198 576642 121488 576716
rect 100896 575058 121488 576642
rect 40404 565351 40428 565352
rect 40404 563045 40405 565351
rect 40404 563044 40428 563045
rect 40138 561975 42446 561976
rect 40138 559669 40139 561975
rect 42445 559669 42446 561975
rect 40138 559668 42446 559669
rect 100896 554084 102480 575058
rect 121184 574906 121488 575058
rect 121198 574864 121488 574906
rect 123240 574864 123530 576716
rect 185798 576882 188130 577128
rect 185798 576656 186088 576882
rect 185784 576483 186088 576656
rect 121198 574584 123530 574864
rect 170937 575030 186088 576483
rect 187840 575030 188130 576882
rect 170937 574921 188130 575030
rect 121198 572784 123530 573030
rect 121198 572728 121488 572784
rect 106766 571144 121488 572728
rect 100860 553626 103852 554084
rect 100860 551460 101430 553626
rect 103522 551460 103852 553626
rect 100860 550972 103852 551460
rect 100896 545334 102480 550972
rect 106766 549804 108350 571144
rect 121184 570974 121488 571144
rect 121198 570932 121488 570974
rect 123240 570932 123530 572784
rect 121198 570652 123530 570932
rect 121198 568942 123530 569188
rect 121198 568716 121488 568942
rect 121184 568610 121488 568716
rect 111760 567090 121488 568610
rect 123240 567090 123530 568942
rect 111760 567026 123530 567090
rect 106354 549502 109178 549804
rect 106354 547336 106858 549502
rect 108950 547336 109178 549502
rect 106354 547098 109178 547336
rect 93214 543750 102480 545334
rect 106766 498256 108350 547098
rect 93214 496672 108350 498256
rect 111760 545514 113344 567026
rect 121198 566810 123530 567026
rect 114747 563203 117455 563204
rect 114747 560497 114748 563203
rect 117454 560497 119479 563203
rect 114747 560496 119479 560497
rect 111760 545174 115256 545514
rect 111760 542488 112142 545174
rect 114828 542488 115256 545174
rect 111760 541920 115256 542488
rect 103002 494539 104586 496672
rect 103002 492957 103003 494539
rect 104585 492957 104586 494539
rect 103002 492956 104586 492957
rect 111760 483970 113344 541920
rect 116773 496039 119479 560496
rect 121184 556994 123516 557240
rect 121184 556768 121474 556994
rect 121170 555184 121474 556768
rect 121184 555142 121474 555184
rect 123226 555142 123516 556994
rect 121184 554862 123516 555142
rect 121198 553450 123530 553696
rect 121198 553224 121488 553450
rect 121184 551640 121488 553224
rect 121198 551598 121488 551640
rect 123240 551598 123530 553450
rect 170937 553119 172499 574921
rect 185798 574750 188130 574921
rect 185798 573242 188130 573488
rect 185798 573016 186088 573242
rect 185784 572929 186088 573016
rect 121198 551318 123530 551598
rect 164479 551557 172499 553119
rect 175957 571390 186088 572929
rect 187840 571390 188130 573242
rect 175957 571367 188130 571390
rect 121198 549846 123530 550092
rect 121198 549620 121488 549846
rect 121184 548036 121488 549620
rect 121198 547994 121488 548036
rect 123240 547994 123530 549846
rect 121198 547714 123530 547994
rect 164479 549156 166041 551557
rect 164479 547596 164480 549156
rect 166040 547596 166041 549156
rect 121198 545914 123530 546160
rect 121198 545688 121488 545914
rect 121184 544104 121488 545688
rect 121198 544062 121488 544104
rect 123240 544062 123530 545914
rect 164479 545521 166041 547596
rect 121198 543782 123530 544062
rect 157613 543959 166041 545521
rect 175957 545187 177519 571367
rect 185798 571110 188130 571367
rect 185798 553434 188130 553680
rect 185798 553208 186088 553434
rect 185784 551624 186088 553208
rect 185798 551582 186088 551624
rect 187840 551582 188130 553434
rect 185798 551302 188130 551582
rect 185798 549390 188130 549636
rect 185798 549164 186088 549390
rect 185784 547580 186088 549164
rect 185798 547538 186088 547580
rect 187840 547538 188130 549390
rect 185798 547258 188130 547538
rect 185798 545752 188130 545998
rect 448623 545981 458103 584769
rect 185798 545526 186088 545752
rect 185784 545187 186088 545526
rect 175957 543900 186088 545187
rect 187840 545187 188130 545752
rect 187840 543900 188373 545187
rect 175957 543625 188373 543900
rect 175957 524271 177519 543625
rect 185798 543620 188130 543625
rect 221885 542099 458480 545981
rect 171643 522709 177519 524271
rect 171643 497921 173205 522709
rect 157885 496359 173205 497921
rect 116773 495450 123695 496039
rect 116773 493598 121488 495450
rect 123240 493598 123695 495450
rect 157885 495437 159447 496359
rect 116773 493333 123695 493598
rect 121198 493318 123530 493333
rect 121198 491518 123530 491764
rect 121198 491292 121488 491518
rect 121184 489708 121488 491292
rect 121198 489666 121488 489708
rect 123240 489666 123530 491518
rect 121198 489386 123530 489666
rect 121198 487914 123530 488160
rect 121198 487688 121488 487914
rect 121184 486104 121488 487688
rect 121198 486062 121488 486104
rect 123240 486062 123530 487914
rect 121198 485782 123530 486062
rect 121170 484326 123502 484572
rect 121170 484100 121460 484326
rect 121156 483970 121460 484100
rect 111760 482474 121460 483970
rect 123212 483970 123502 484326
rect 123212 482474 123514 483970
rect 111760 482386 123514 482474
rect 33508 480757 35816 480758
rect 33508 478451 33509 480757
rect 35815 478451 35816 480757
rect 33508 478450 35816 478451
rect 29694 477029 32002 477030
rect 29694 474723 29695 477029
rect 32001 474723 32002 477029
rect 29694 474722 32002 474723
rect 111760 461048 113344 482386
rect 121170 482194 123502 482386
rect 93156 459464 113344 461048
<< via4 >>
rect 40428 565351 42736 565352
rect 40428 563045 42711 565351
rect 42711 563045 42736 565351
rect 40428 563044 42736 563045
rect 40162 559692 42422 561952
rect 487752 566680 503872 566681
rect 487752 550562 487753 566680
rect 487753 550562 503871 566680
rect 503871 550562 503872 566680
rect 487752 550561 503872 550562
rect 33532 478474 35792 480734
rect 29718 474746 31978 477006
rect 527393 481837 543845 481838
rect 527393 465387 527394 481837
rect 527394 465387 543844 481837
rect 543844 465387 543845 481837
rect 527393 465386 543845 465387
<< metal5 >>
rect 99272 605640 194538 607948
rect 225312 605640 260148 607948
rect 252960 567500 260148 605640
rect 252960 566681 513241 567500
rect 40404 565352 42760 565376
rect 40404 563044 40428 565352
rect 42736 563044 64980 565352
rect 96858 563044 127852 565352
rect 159520 563044 195514 565352
rect 40404 563020 42760 563044
rect 40138 561952 64596 561976
rect 40138 559692 40162 561952
rect 42422 559692 64596 561952
rect 40138 559668 64596 559692
rect 96858 559668 130612 561976
rect 162222 559668 197526 561976
rect 252960 550561 487752 566681
rect 503872 550561 513241 566681
rect 252960 546234 513241 550561
rect 98838 520694 127800 523002
rect 252960 521196 260148 546234
rect 252960 519380 260568 521196
rect 96728 517072 128926 519380
rect 162038 519269 195206 519380
rect 162038 517072 196477 519269
rect 223220 518888 260568 519380
rect 223220 517072 260148 518888
rect 189832 487858 196477 517072
rect 252960 516960 255268 517072
rect 257840 515886 260148 517072
rect 189832 481838 544282 487858
rect 33508 480734 65058 480758
rect 33508 478474 33532 480734
rect 35792 478474 65058 480734
rect 33508 478450 65058 478474
rect 29694 477006 64134 477030
rect 29694 474746 29718 477006
rect 31978 474746 64134 477006
rect 29694 474722 64134 474746
rect 95552 474722 136672 477030
rect 189832 465386 527393 481838
rect 543845 465386 544282 481838
rect 189832 464706 544282 465386
rect 189832 434786 196477 464706
rect 95624 432478 196477 434786
rect 191278 432148 193586 432478
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use analog_neuron  analog_neuron_3 ~/Documents/AnalogNeuron/opamp
timestamp 1624077225
transform 1 0 43138 0 -1 895902
box 18328 415144 58222 463464
use analog_neuron  analog_neuron_1
array 0 2 64338 0 0 48320
timestamp 1624077225
transform 1 0 43294 0 -1 980496
box 18328 415144 58222 463464
use analog_neuron  analog_neuron_4
array 0 1 64628 0 0 -47922
timestamp 1624077225
transform 1 0 43154 0 1 59578
box 18328 415144 58222 463464
use analog_neuron  analog_neuron_0
array 0 2 64338 0 0 48320
timestamp 1624077225
transform 1 0 43310 0 1 144524
box 18328 415144 58222 463464
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
rlabel poly 130634 568376 130638 568406 7 p2
port 2 w
rlabel polycont 129954 568376 129958 568406 3 p1
port 1 e
rlabel poly 130604 556316 130608 556346 7 p2
port 2 w
rlabel polycont 129924 556316 129928 556346 3 p1
port 1 e
rlabel poly 130740 483684 130744 483714 7 p2
port 2 w
rlabel polycont 130060 483684 130064 483714 3 p1
port 1 e
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
