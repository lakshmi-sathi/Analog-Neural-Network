magic
tech sky130A
magscale 1 2
timestamp 1627923075
<< xpolycontact >>
rect -35 638 35 1070
rect -35 -1070 35 -638
<< xpolyres >>
rect -35 -638 35 638
<< viali >>
rect -19 655 19 1052
rect -19 -1052 19 -655
<< metal1 >>
rect -25 1052 25 1064
rect -25 655 -19 1052
rect 19 655 25 1052
rect -25 643 25 655
rect -25 -655 25 -643
rect -25 -1052 -19 -655
rect 19 -1052 25 -655
rect -25 -1064 25 -1052
<< res0p35 >>
rect -37 -640 37 640
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 6.38 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 37.142k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
