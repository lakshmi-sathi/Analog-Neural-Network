magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_s >>
rect -10 228 102 238
rect -10 172 32 228
rect -10 162 102 172
rect 694 84 1052 190
rect 862 22 884 84
rect 958 22 1052 84
rect 826 -2 1052 22
rect -22 -34 100 -26
rect -22 -98 25 -34
rect 826 -40 920 -2
rect 958 -40 1052 -2
rect -22 -104 100 -98
rect 826 -146 1052 -40
rect 862 -147 1052 -146
<< nwell >>
rect 263 52 481 85
rect 263 50 506 52
rect 263 -181 481 50
rect 884 -2 958 84
rect 848 -40 958 -2
rect 856 -146 858 -128
rect 263 -245 537 -181
rect 884 -246 958 -40
<< pwell >>
rect 860 154 942 238
rect 862 -2 884 22
rect 862 -146 884 -40
<< nmos >>
rect 359 157 389 241
<< pmos >>
rect 357 -145 387 23
<< ndiff >>
rect 301 216 359 241
rect 301 182 313 216
rect 347 182 359 216
rect 301 157 359 182
rect 389 216 447 241
rect 389 182 401 216
rect 435 182 447 216
rect 389 157 447 182
rect 854 154 860 238
<< pdiff >>
rect 299 -10 357 23
rect 299 -44 311 -10
rect 345 -44 357 -10
rect 299 -78 357 -44
rect 299 -112 311 -78
rect 345 -112 357 -78
rect 299 -145 357 -112
rect 387 -10 445 23
rect 387 -44 399 -10
rect 433 -44 445 -10
rect 387 -78 445 -44
rect 387 -112 399 -78
rect 433 -112 445 -78
rect 387 -145 445 -112
rect 856 -146 862 22
<< ndiffc >>
rect 313 182 347 216
rect 401 182 435 216
<< pdiffc >>
rect 311 -44 345 -10
rect 311 -112 345 -78
rect 399 -44 433 -10
rect 399 -112 433 -78
<< psubdiff >>
rect 860 213 942 238
rect 860 179 884 213
rect 918 179 942 213
rect 860 154 942 179
<< nsubdiff >>
rect 862 -48 920 22
rect 862 -82 884 -48
rect 918 -82 920 -48
rect 862 -146 920 -82
<< psubdiffcont >>
rect 884 179 918 213
<< nsubdiffcont >>
rect 884 -82 918 -48
<< poly >>
rect 341 313 407 329
rect 341 279 357 313
rect 391 279 407 313
rect 341 263 407 279
rect 359 241 389 263
rect 359 131 389 157
rect 357 23 387 49
rect 770 35 800 154
rect 357 -176 387 -145
rect 339 -192 405 -176
rect 339 -226 355 -192
rect 389 -226 405 -192
rect 339 -242 405 -226
<< polycont >>
rect 357 279 391 313
rect 355 -226 389 -192
<< locali >>
rect 156 331 393 373
rect 156 -120 198 331
rect 341 313 393 331
rect 540 356 714 398
rect 341 279 357 313
rect 391 279 407 313
rect 540 298 608 356
rect 540 292 582 298
rect 313 216 347 245
rect 401 217 435 245
rect 678 242 714 356
rect 678 234 754 242
rect 311 182 313 209
rect 311 -8 347 182
rect 345 -44 347 -8
rect 311 -78 347 -44
rect 345 -114 347 -78
rect 156 -191 200 -120
rect 311 -135 347 -114
rect 397 216 435 217
rect 397 182 401 216
rect 397 153 435 182
rect 397 -8 433 153
rect 397 -44 399 -8
rect 397 -78 433 -44
rect 397 -114 399 -78
rect 397 -127 433 -114
rect 311 -149 345 -135
rect 399 -149 433 -127
rect 511 -135 547 209
rect 597 -127 633 217
rect 678 152 758 234
rect 884 213 918 246
rect 884 148 918 179
rect 882 -48 920 2
rect 882 -82 884 -48
rect 882 -130 920 -82
rect 156 -233 204 -191
rect 338 -192 406 -190
rect 338 -226 355 -192
rect 389 -226 406 -192
rect 542 -226 780 -192
rect 156 -304 200 -233
rect 338 -234 406 -226
rect 642 -304 686 -226
rect 156 -348 686 -304
<< viali >>
rect 357 279 391 313
rect 313 182 347 216
rect 311 -10 345 -8
rect 311 -42 345 -10
rect 311 -112 345 -80
rect 311 -114 345 -112
rect 401 182 435 216
rect 399 -10 433 -8
rect 399 -42 433 -10
rect 399 -112 433 -80
rect 399 -114 433 -112
rect 884 179 918 213
rect 886 -82 918 -48
rect 918 -82 920 -48
rect 355 -226 389 -192
<< metal1 >>
rect 173 367 606 429
rect 173 -181 235 367
rect 340 319 406 326
rect 544 325 606 367
rect 854 390 940 405
rect 854 338 872 390
rect 924 338 940 390
rect 340 313 407 319
rect 340 279 357 313
rect 391 279 407 313
rect 340 270 407 279
rect 543 271 607 325
rect 754 266 814 322
rect 307 240 353 241
rect 284 223 354 240
rect 284 171 291 223
rect 343 216 354 223
rect 347 182 354 216
rect 343 171 354 182
rect 284 154 354 171
rect 395 236 441 241
rect 395 216 458 236
rect 594 223 660 242
rect 854 238 940 338
rect 395 182 401 216
rect 435 182 458 216
rect 395 157 458 182
rect 396 156 458 157
rect 506 124 556 216
rect 594 171 600 223
rect 652 171 660 223
rect 594 154 660 171
rect 474 114 558 124
rect 474 62 489 114
rect 541 62 558 114
rect 474 52 558 62
rect 506 50 558 52
rect 396 23 458 24
rect 305 22 351 23
rect 286 -8 351 22
rect 286 -42 311 -8
rect 345 -42 351 -8
rect 286 -80 351 -42
rect 286 -114 311 -80
rect 345 -114 351 -80
rect 286 -144 351 -114
rect 305 -145 351 -144
rect 393 -8 458 23
rect 506 10 556 50
rect 393 -42 399 -8
rect 433 -35 458 -8
rect 718 -18 762 236
rect 816 213 940 238
rect 816 179 884 213
rect 918 179 940 213
rect 816 164 940 179
rect 848 -30 936 -2
rect 393 -80 406 -42
rect 824 -48 936 -30
rect 824 -50 886 -48
rect 393 -114 399 -80
rect 433 -114 458 -87
rect 393 -145 458 -114
rect 396 -146 458 -145
rect 806 -82 886 -50
rect 920 -82 936 -48
rect 806 -146 936 -82
rect 339 -181 405 -179
rect 173 -192 405 -181
rect 173 -226 355 -192
rect 389 -226 405 -192
rect 173 -243 405 -226
rect 537 -235 601 -185
rect 752 -232 820 -184
rect 862 -206 936 -146
rect 545 -248 596 -235
rect 862 -258 874 -206
rect 926 -258 936 -206
rect 862 -270 936 -258
<< via1 >>
rect 872 338 924 390
rect 291 216 343 223
rect 291 182 313 216
rect 313 182 343 216
rect 291 171 343 182
rect 600 171 652 223
rect 489 62 541 114
rect 406 -42 433 -35
rect 433 -42 458 -35
rect 406 -80 458 -42
rect 406 -87 433 -80
rect 433 -87 458 -80
rect 874 -258 926 -206
<< metal2 >>
rect 858 390 938 402
rect 858 338 872 390
rect 924 338 938 390
rect 858 324 938 338
rect 594 240 660 242
rect 594 238 978 240
rect 20 228 350 238
rect 20 172 32 228
rect 88 223 350 228
rect 88 172 291 223
rect 20 171 291 172
rect 343 171 350 223
rect 20 158 350 171
rect 594 223 996 238
rect 594 171 600 223
rect 652 171 996 223
rect 594 154 996 171
rect 484 116 546 126
rect 484 60 487 116
rect 543 60 546 116
rect 484 50 546 60
rect 926 104 996 154
rect 926 30 1124 104
rect 22 -38 92 -22
rect 926 -24 996 30
rect 22 -94 29 -38
rect 85 -94 92 -38
rect 22 -110 92 -94
rect 400 -35 996 -24
rect 400 -87 406 -35
rect 458 -87 996 -35
rect 400 -98 996 -87
rect 654 -100 996 -98
rect 926 -102 996 -100
rect 866 -206 936 -198
rect 866 -258 874 -206
rect 926 -258 936 -206
rect 866 -268 936 -258
<< via2 >>
rect 32 172 88 228
rect 487 114 543 116
rect 487 62 489 114
rect 489 62 541 114
rect 541 62 543 114
rect 487 60 543 62
rect 29 -94 85 -38
<< metal3 >>
rect -10 228 102 238
rect -10 172 32 228
rect 88 172 102 228
rect -10 162 102 172
rect 468 116 558 138
rect 468 98 487 116
rect 466 78 487 98
rect 4 60 487 78
rect 543 60 558 116
rect 4 26 558 60
rect 4 18 544 26
rect 8 -34 110 18
rect 8 -98 25 -34
rect 89 -98 110 -34
rect 8 -114 110 -98
<< via3 >>
rect 25 -38 89 -34
rect 25 -94 29 -38
rect 29 -94 85 -38
rect 85 -94 89 -38
rect 25 -98 89 -94
<< metal4 >>
rect -22 -34 100 -26
rect -22 -98 25 -34
rect 89 -98 100 -34
rect -22 -104 100 -98
use sky130_fd_pr__pfet_01v8_EMKQNQ  sky130_fd_pr__pfet_01v8_EMKQNQ_0
timestamp 1627926120
transform 1 0 785 0 1 -98
box -109 -148 267 288
use sky130_fd_pr__nfet_01v8_SLJCGW  sky130_fd_pr__nfet_01v8_SLJCGW_0
timestamp 1627926120
transform 1 0 574 0 1 230
box -73 -99 73 99
use sky130_fd_pr__nfet_01v8_SLJCGW  sky130_fd_pr__nfet_01v8_SLJCGW_1
timestamp 1627926120
transform 1 0 785 0 1 227
box -73 -99 73 99
use sky130_fd_pr__pfet_01v8_E6WEYA  sky130_fd_pr__pfet_01v8_E6WEYA_0
timestamp 1627926120
transform -1 0 572 0 -1 -97
box -109 -182 109 148
<< labels >>
rlabel locali s 160 -340 192 -134 4 sel
port 1 nsew
rlabel metal2 s 860 326 936 400 4 GND
port 2 nsew
rlabel metal2 s 868 -266 932 -200 4 VDD
port 3 nsew
rlabel metal3 s 0 168 98 234 4 in1
port 4 nsew
rlabel metal4 s -16 -102 98 -28 4 in2
port 5 nsew
rlabel metal2 s 948 36 1116 98 4 out
port 6 nsew
<< end >>
