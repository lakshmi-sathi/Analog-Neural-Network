magic
tech sky130A
magscale 1 2
timestamp 1627921586
<< xpolycontact >>
rect -35 893 35 1325
rect -35 -1325 35 -893
<< xpolyres >>
rect -35 -893 35 893
<< viali >>
rect -19 910 19 1307
rect -19 -1307 19 -910
<< metal1 >>
rect -25 1307 25 1319
rect -25 910 -19 1307
rect 19 910 25 1307
rect -25 898 25 910
rect -25 -910 25 -898
rect -25 -1307 -19 -910
rect 19 -1307 25 -910
rect -25 -1319 25 -1307
<< res0p35 >>
rect -37 -895 37 895
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 8.93 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 51.714k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
