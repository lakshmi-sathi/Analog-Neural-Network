magic
tech sky130A
magscale 1 2
timestamp 1627111729
<< xpolycontact >>
rect -141 165 141 597
rect -141 -597 141 -165
<< xpolyres >>
rect -141 -165 141 165
<< viali >>
rect -125 182 125 579
rect -125 -579 125 -182
<< metal1 >>
rect -131 579 131 591
rect -131 182 -125 579
rect 125 182 131 579
rect -131 170 131 182
rect -131 -182 131 -170
rect -131 -579 -125 -182
rect 125 -579 131 -182
rect -131 -591 131 -579
<< res1p41 >>
rect -143 -167 143 167
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string parameters w 1.410 l 1.65 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 2.51k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
