magic
tech sky130A
magscale 1 2
timestamp 1627800883
<< poly >>
rect 3963 675 4060 701
rect 3967 671 4060 675
rect 4030 623 4060 671
<< locali >>
rect 50 -128 4114 -118
rect 50 -206 62 -128
rect 4102 -206 4114 -128
rect 50 -216 4114 -206
<< viali >>
rect 62 -206 4102 -128
<< metal1 >>
rect 76 654 3980 706
rect 126 620 188 622
rect 318 620 380 622
rect 510 620 572 622
rect 702 620 764 622
rect 894 620 956 622
rect 1086 620 1148 622
rect 1278 620 1340 622
rect 1470 620 1532 622
rect 1662 620 1724 622
rect 1854 620 1916 622
rect 2046 620 2108 622
rect 2238 620 2300 622
rect 2430 620 2492 622
rect 2622 620 2684 622
rect 2814 620 2876 622
rect 3006 620 3068 622
rect 3198 620 3260 622
rect 3390 620 3452 622
rect 3582 620 3644 622
rect 3774 620 3836 622
rect 3966 620 4028 622
rect 126 614 190 620
rect 126 364 132 614
rect 184 364 190 614
rect 318 614 382 620
rect 318 364 324 614
rect 376 364 382 614
rect 510 614 574 620
rect 510 364 516 614
rect 568 364 574 614
rect 702 614 766 620
rect 702 364 708 614
rect 760 364 766 614
rect 894 614 958 620
rect 894 364 900 614
rect 952 364 958 614
rect 1086 614 1150 620
rect 1086 364 1092 614
rect 1144 364 1150 614
rect 1278 614 1342 620
rect 1278 364 1284 614
rect 1336 364 1342 614
rect 1470 614 1534 620
rect 1470 364 1476 614
rect 1528 364 1534 614
rect 1662 614 1726 620
rect 1662 364 1668 614
rect 1720 364 1726 614
rect 1854 614 1918 620
rect 1854 364 1860 614
rect 1912 364 1918 614
rect 2046 614 2110 620
rect 2046 364 2052 614
rect 2104 364 2110 614
rect 2238 614 2302 620
rect 2238 364 2244 614
rect 2296 364 2302 614
rect 2430 614 2494 620
rect 2430 364 2436 614
rect 2488 364 2494 614
rect 2622 614 2686 620
rect 2622 364 2628 614
rect 2680 364 2686 614
rect 2814 614 2878 620
rect 2814 364 2820 614
rect 2872 364 2878 614
rect 3006 614 3070 620
rect 3006 364 3012 614
rect 3064 364 3070 614
rect 3198 614 3262 620
rect 3198 364 3204 614
rect 3256 364 3262 614
rect 3390 614 3454 620
rect 3390 364 3396 614
rect 3448 364 3454 614
rect 3582 614 3646 620
rect 3582 364 3588 614
rect 3640 364 3646 614
rect 3774 614 3838 620
rect 3774 364 3780 614
rect 3832 364 3838 614
rect 3966 614 4030 620
rect 3966 364 3972 614
rect 4024 364 4030 614
rect 30 30 36 284
rect 88 30 94 284
rect 30 24 94 30
rect 222 30 228 284
rect 280 30 286 284
rect 222 24 286 30
rect 414 30 420 284
rect 472 30 478 284
rect 414 24 478 30
rect 606 30 612 284
rect 664 30 670 284
rect 606 24 670 30
rect 798 30 804 284
rect 856 30 862 284
rect 798 24 862 30
rect 990 30 996 284
rect 1048 30 1054 284
rect 990 24 1054 30
rect 1182 30 1188 284
rect 1240 30 1246 284
rect 1182 24 1246 30
rect 1374 30 1380 284
rect 1432 30 1438 284
rect 1374 24 1438 30
rect 1566 30 1572 284
rect 1624 30 1630 284
rect 1566 24 1630 30
rect 1758 30 1764 284
rect 1816 30 1822 284
rect 1758 24 1822 30
rect 1950 30 1956 284
rect 2008 30 2014 284
rect 1950 24 2014 30
rect 2142 30 2148 284
rect 2200 30 2206 284
rect 2142 24 2206 30
rect 2334 30 2340 284
rect 2392 30 2398 284
rect 2334 24 2398 30
rect 2526 30 2532 284
rect 2584 30 2590 284
rect 2526 24 2590 30
rect 2718 30 2724 284
rect 2776 30 2782 284
rect 2718 24 2782 30
rect 2910 30 2916 284
rect 2968 30 2974 284
rect 2910 24 2974 30
rect 3102 30 3108 284
rect 3160 30 3166 284
rect 3102 24 3166 30
rect 3294 30 3300 284
rect 3352 30 3358 284
rect 3294 24 3358 30
rect 3486 30 3492 284
rect 3544 30 3550 284
rect 3486 24 3550 30
rect 3678 30 3684 284
rect 3736 30 3742 284
rect 3678 24 3742 30
rect 3870 30 3876 284
rect 3928 30 3934 284
rect 3870 24 3934 30
rect 4062 30 4068 284
rect 4120 30 4126 284
rect 4062 24 4126 30
rect 172 -60 4076 -8
rect 50 -128 4114 -116
rect 50 -208 62 -128
rect 4104 -208 4114 -128
rect 50 -220 4114 -208
<< via1 >>
rect 132 364 184 614
rect 324 364 376 614
rect 516 364 568 614
rect 708 364 760 614
rect 900 364 952 614
rect 1092 364 1144 614
rect 1284 364 1336 614
rect 1476 364 1528 614
rect 1668 364 1720 614
rect 1860 364 1912 614
rect 2052 364 2104 614
rect 2244 364 2296 614
rect 2436 364 2488 614
rect 2628 364 2680 614
rect 2820 364 2872 614
rect 3012 364 3064 614
rect 3204 364 3256 614
rect 3396 364 3448 614
rect 3588 364 3640 614
rect 3780 364 3832 614
rect 3972 364 4024 614
rect 36 30 88 284
rect 228 30 280 284
rect 420 30 472 284
rect 612 30 664 284
rect 804 30 856 284
rect 996 30 1048 284
rect 1188 30 1240 284
rect 1380 30 1432 284
rect 1572 30 1624 284
rect 1764 30 1816 284
rect 1956 30 2008 284
rect 2148 30 2200 284
rect 2340 30 2392 284
rect 2532 30 2584 284
rect 2724 30 2776 284
rect 2916 30 2968 284
rect 3108 30 3160 284
rect 3300 30 3352 284
rect 3492 30 3544 284
rect 3684 30 3736 284
rect 3876 30 3928 284
rect 4068 30 4120 284
rect 62 -206 4102 -128
rect 4102 -206 4104 -128
rect 62 -208 4104 -206
<< metal2 >>
rect 126 620 188 622
rect 318 620 380 622
rect 510 620 572 622
rect 702 620 764 622
rect 894 620 956 622
rect 1086 620 1148 622
rect 1278 620 1340 622
rect 1470 620 1532 622
rect 1662 620 1724 622
rect 1854 620 1916 622
rect 2046 620 2108 622
rect 2238 620 2300 622
rect 2430 620 2492 622
rect 2622 620 2684 622
rect 2814 620 2876 622
rect 3006 620 3068 622
rect 3198 620 3260 622
rect 3390 620 3452 622
rect 3582 620 3644 622
rect 3774 620 3836 622
rect 3966 620 4028 622
rect 126 614 190 620
rect 126 612 132 614
rect 184 612 190 614
rect 126 364 130 612
rect 186 364 190 612
rect 126 354 190 364
rect 318 614 382 620
rect 318 612 324 614
rect 376 612 382 614
rect 318 364 322 612
rect 378 364 382 612
rect 318 354 382 364
rect 510 614 574 620
rect 510 612 516 614
rect 568 612 574 614
rect 510 364 514 612
rect 570 364 574 612
rect 510 354 574 364
rect 702 614 766 620
rect 702 612 708 614
rect 760 612 766 614
rect 702 364 706 612
rect 762 364 766 612
rect 702 354 766 364
rect 894 614 958 620
rect 894 612 900 614
rect 952 612 958 614
rect 894 364 898 612
rect 954 364 958 612
rect 894 354 958 364
rect 1086 614 1150 620
rect 1086 612 1092 614
rect 1144 612 1150 614
rect 1086 364 1090 612
rect 1146 364 1150 612
rect 1086 354 1150 364
rect 1278 614 1342 620
rect 1278 612 1284 614
rect 1336 612 1342 614
rect 1278 364 1282 612
rect 1338 364 1342 612
rect 1278 354 1342 364
rect 1470 614 1534 620
rect 1470 612 1476 614
rect 1528 612 1534 614
rect 1470 364 1474 612
rect 1530 364 1534 612
rect 1470 354 1534 364
rect 1662 614 1726 620
rect 1662 612 1668 614
rect 1720 612 1726 614
rect 1662 364 1666 612
rect 1722 364 1726 612
rect 1662 354 1726 364
rect 1854 614 1918 620
rect 1854 612 1860 614
rect 1912 612 1918 614
rect 1854 364 1858 612
rect 1914 364 1918 612
rect 1854 354 1918 364
rect 2046 614 2110 620
rect 2046 612 2052 614
rect 2104 612 2110 614
rect 2046 364 2050 612
rect 2106 364 2110 612
rect 2046 354 2110 364
rect 2238 614 2302 620
rect 2238 612 2244 614
rect 2296 612 2302 614
rect 2238 364 2242 612
rect 2298 364 2302 612
rect 2238 354 2302 364
rect 2430 614 2494 620
rect 2430 612 2436 614
rect 2488 612 2494 614
rect 2430 364 2434 612
rect 2490 364 2494 612
rect 2430 354 2494 364
rect 2622 614 2686 620
rect 2622 612 2628 614
rect 2680 612 2686 614
rect 2622 364 2626 612
rect 2682 364 2686 612
rect 2622 354 2686 364
rect 2814 614 2878 620
rect 2814 612 2820 614
rect 2872 612 2878 614
rect 2814 364 2818 612
rect 2874 364 2878 612
rect 2814 354 2878 364
rect 3006 614 3070 620
rect 3006 612 3012 614
rect 3064 612 3070 614
rect 3006 364 3010 612
rect 3066 364 3070 612
rect 3006 354 3070 364
rect 3198 614 3262 620
rect 3198 612 3204 614
rect 3256 612 3262 614
rect 3198 364 3202 612
rect 3258 364 3262 612
rect 3198 354 3262 364
rect 3390 614 3454 620
rect 3390 612 3396 614
rect 3448 612 3454 614
rect 3390 364 3394 612
rect 3450 364 3454 612
rect 3390 354 3454 364
rect 3582 614 3646 620
rect 3582 612 3588 614
rect 3640 612 3646 614
rect 3582 364 3586 612
rect 3642 364 3646 612
rect 3582 354 3646 364
rect 3774 614 3838 620
rect 3774 612 3780 614
rect 3832 612 3838 614
rect 3774 364 3778 612
rect 3834 364 3838 612
rect 3774 354 3838 364
rect 3966 614 4030 620
rect 3966 612 3972 614
rect 4024 612 4030 614
rect 3966 364 3970 612
rect 4026 364 4030 612
rect 3966 354 4030 364
rect 30 30 36 284
rect 88 30 94 284
rect 30 -76 94 30
rect 222 30 228 284
rect 280 30 286 284
rect 222 -76 286 30
rect 414 30 420 284
rect 472 30 478 284
rect 414 -76 478 30
rect 606 30 612 284
rect 664 30 670 284
rect 606 -76 670 30
rect 798 30 804 284
rect 856 30 862 284
rect 798 -76 862 30
rect 990 30 996 284
rect 1048 30 1054 284
rect 990 -76 1054 30
rect 1182 30 1188 284
rect 1240 30 1246 284
rect 1182 -76 1246 30
rect 1374 30 1380 284
rect 1432 30 1438 284
rect 1374 -76 1438 30
rect 1566 30 1572 284
rect 1624 30 1630 284
rect 1566 -76 1630 30
rect 1758 30 1764 284
rect 1816 30 1822 284
rect 1758 -76 1822 30
rect 1950 30 1956 284
rect 2008 30 2014 284
rect 1950 -76 2014 30
rect 2142 30 2148 284
rect 2200 30 2206 284
rect 2142 -76 2206 30
rect 2334 30 2340 284
rect 2392 30 2398 284
rect 2334 -76 2398 30
rect 2526 30 2532 284
rect 2584 30 2590 284
rect 2526 -76 2590 30
rect 2718 30 2724 284
rect 2776 30 2782 284
rect 2718 -76 2782 30
rect 2910 30 2916 284
rect 2968 30 2974 284
rect 2910 -76 2974 30
rect 3102 30 3108 284
rect 3160 30 3166 284
rect 3102 -76 3166 30
rect 3294 30 3300 284
rect 3352 30 3358 284
rect 3294 -76 3358 30
rect 3486 30 3492 284
rect 3544 30 3550 284
rect 3486 -76 3550 30
rect 3678 30 3684 284
rect 3736 30 3742 284
rect 3678 -76 3742 30
rect 3870 30 3876 284
rect 3928 30 3934 284
rect 3870 -76 3934 30
rect 4062 30 4068 284
rect 4120 30 4126 284
rect 4062 -76 4126 30
rect 24 -128 4130 -76
rect 24 -208 62 -128
rect 4104 -208 4130 -128
rect 24 -284 4130 -208
rect 24 -320 4128 -284
<< via2 >>
rect 130 364 132 612
rect 132 364 184 612
rect 184 364 186 612
rect 322 364 324 612
rect 324 364 376 612
rect 376 364 378 612
rect 514 364 516 612
rect 516 364 568 612
rect 568 364 570 612
rect 706 364 708 612
rect 708 364 760 612
rect 760 364 762 612
rect 898 364 900 612
rect 900 364 952 612
rect 952 364 954 612
rect 1090 364 1092 612
rect 1092 364 1144 612
rect 1144 364 1146 612
rect 1282 364 1284 612
rect 1284 364 1336 612
rect 1336 364 1338 612
rect 1474 364 1476 612
rect 1476 364 1528 612
rect 1528 364 1530 612
rect 1666 364 1668 612
rect 1668 364 1720 612
rect 1720 364 1722 612
rect 1858 364 1860 612
rect 1860 364 1912 612
rect 1912 364 1914 612
rect 2050 364 2052 612
rect 2052 364 2104 612
rect 2104 364 2106 612
rect 2242 364 2244 612
rect 2244 364 2296 612
rect 2296 364 2298 612
rect 2434 364 2436 612
rect 2436 364 2488 612
rect 2488 364 2490 612
rect 2626 364 2628 612
rect 2628 364 2680 612
rect 2680 364 2682 612
rect 2818 364 2820 612
rect 2820 364 2872 612
rect 2872 364 2874 612
rect 3010 364 3012 612
rect 3012 364 3064 612
rect 3064 364 3066 612
rect 3202 364 3204 612
rect 3204 364 3256 612
rect 3256 364 3258 612
rect 3394 364 3396 612
rect 3396 364 3448 612
rect 3448 364 3450 612
rect 3586 364 3588 612
rect 3588 364 3640 612
rect 3640 364 3642 612
rect 3778 364 3780 612
rect 3780 364 3832 612
rect 3832 364 3834 612
rect 3970 364 3972 612
rect 3972 364 4024 612
rect 4024 364 4026 612
<< metal3 >>
rect 124 728 4032 814
rect 124 612 192 728
rect 124 364 130 612
rect 186 364 192 612
rect 124 354 192 364
rect 316 612 384 728
rect 316 364 322 612
rect 378 364 384 612
rect 316 354 384 364
rect 508 612 576 728
rect 508 364 514 612
rect 570 364 576 612
rect 508 354 576 364
rect 700 612 768 728
rect 700 364 706 612
rect 762 364 768 612
rect 700 354 768 364
rect 892 612 960 728
rect 892 364 898 612
rect 954 364 960 612
rect 892 354 960 364
rect 1084 612 1152 728
rect 1084 364 1090 612
rect 1146 364 1152 612
rect 1084 354 1152 364
rect 1276 612 1344 728
rect 1276 364 1282 612
rect 1338 364 1344 612
rect 1276 354 1344 364
rect 1468 612 1536 728
rect 1468 364 1474 612
rect 1530 364 1536 612
rect 1468 354 1536 364
rect 1660 612 1728 728
rect 1660 364 1666 612
rect 1722 364 1728 612
rect 1660 354 1728 364
rect 1852 612 1920 728
rect 1852 364 1858 612
rect 1914 364 1920 612
rect 1852 354 1920 364
rect 2044 612 2112 728
rect 2044 364 2050 612
rect 2106 364 2112 612
rect 2044 354 2112 364
rect 2236 612 2304 728
rect 2236 364 2242 612
rect 2298 364 2304 612
rect 2236 354 2304 364
rect 2428 612 2496 728
rect 2428 364 2434 612
rect 2490 364 2496 612
rect 2428 354 2496 364
rect 2620 612 2688 728
rect 2620 364 2626 612
rect 2682 364 2688 612
rect 2620 354 2688 364
rect 2812 612 2880 728
rect 2812 364 2818 612
rect 2874 364 2880 612
rect 2812 354 2880 364
rect 3004 612 3072 728
rect 3004 364 3010 612
rect 3066 364 3072 612
rect 3004 354 3072 364
rect 3196 612 3264 728
rect 3196 364 3202 612
rect 3258 364 3264 612
rect 3196 354 3264 364
rect 3388 612 3456 728
rect 3388 364 3394 612
rect 3450 364 3456 612
rect 3388 354 3456 364
rect 3580 612 3648 728
rect 3580 364 3586 612
rect 3642 364 3648 612
rect 3580 354 3648 364
rect 3772 612 3840 728
rect 3772 364 3778 612
rect 3834 364 3840 612
rect 3772 354 3840 364
rect 3964 612 4032 728
rect 3964 364 3970 612
rect 4026 364 4032 612
rect 3964 354 4032 364
use sky130_fd_pr__nfet_01v8_4PXCG5  sky130_fd_pr__nfet_01v8_4PXCG5_0
timestamp 1627727346
transform 1 0 2077 0 -1 323
box -2183 -510 2183 510
<< labels >>
rlabel metal2 28 -318 4124 -206 1 GND
port 2 n
rlabel metal1 80 656 3976 704 1 gate
port 4 n
rlabel metal3 124 748 4024 810 1 vl
port 5 n
<< end >>
