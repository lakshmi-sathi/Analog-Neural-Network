magic
tech sky130A
magscale 1 2
timestamp 1628027270
<< xpolycontact >>
rect -35 234 35 666
rect -35 -666 35 -234
<< xpolyres >>
rect -35 -234 35 234
<< viali >>
rect -19 251 19 648
rect -19 -648 19 -251
<< metal1 >>
rect -25 648 25 660
rect -25 251 -19 648
rect 19 251 25 648
rect -25 239 25 251
rect -25 -251 25 -239
rect -25 -648 -19 -251
rect 19 -648 25 -251
rect -25 -660 25 -648
<< res0p35 >>
rect -37 -236 37 236
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 2.34 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 14.057k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
