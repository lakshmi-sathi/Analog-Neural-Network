magic
tech sky130A
magscale 1 2
timestamp 1626793425
<< error_p >>
rect -845 641 -787 647
rect -653 641 -595 647
rect -461 641 -403 647
rect -269 641 -211 647
rect -77 641 -19 647
rect 115 641 173 647
rect 307 641 365 647
rect 499 641 557 647
rect 691 641 749 647
rect -845 607 -833 641
rect -653 607 -641 641
rect -461 607 -449 641
rect -269 607 -257 641
rect -77 607 -65 641
rect 115 607 127 641
rect 307 607 319 641
rect 499 607 511 641
rect 691 607 703 641
rect -845 601 -787 607
rect -653 601 -595 607
rect -461 601 -403 607
rect -269 601 -211 607
rect -77 601 -19 607
rect 115 601 173 607
rect 307 601 365 607
rect 499 601 557 607
rect 691 601 749 607
rect -749 71 -691 77
rect -557 71 -499 77
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect 595 71 653 77
rect 787 71 845 77
rect -749 37 -737 71
rect -557 37 -545 71
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect 595 37 607 71
rect 787 37 799 71
rect -749 31 -691 37
rect -557 31 -499 37
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect 595 31 653 37
rect 787 31 845 37
rect -749 -37 -691 -31
rect -557 -37 -499 -31
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect 595 -37 653 -31
rect 787 -37 845 -31
rect -749 -71 -737 -37
rect -557 -71 -545 -37
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect 595 -71 607 -37
rect 787 -71 799 -37
rect -749 -77 -691 -71
rect -557 -77 -499 -71
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect 595 -77 653 -71
rect 787 -77 845 -71
rect -845 -607 -787 -601
rect -653 -607 -595 -601
rect -461 -607 -403 -601
rect -269 -607 -211 -601
rect -77 -607 -19 -601
rect 115 -607 173 -601
rect 307 -607 365 -601
rect 499 -607 557 -601
rect 691 -607 749 -601
rect -845 -641 -833 -607
rect -653 -641 -641 -607
rect -461 -641 -449 -607
rect -269 -641 -257 -607
rect -77 -641 -65 -607
rect 115 -641 127 -607
rect 307 -641 319 -607
rect 499 -641 511 -607
rect 691 -641 703 -607
rect -845 -647 -787 -641
rect -653 -647 -595 -641
rect -461 -647 -403 -641
rect -269 -647 -211 -641
rect -77 -647 -19 -641
rect 115 -647 173 -641
rect 307 -647 365 -641
rect 499 -647 557 -641
rect 691 -647 749 -641
<< nwell >>
rect -1031 -779 1031 779
<< pmos >>
rect -831 118 -801 560
rect -735 118 -705 560
rect -639 118 -609 560
rect -543 118 -513 560
rect -447 118 -417 560
rect -351 118 -321 560
rect -255 118 -225 560
rect -159 118 -129 560
rect -63 118 -33 560
rect 33 118 63 560
rect 129 118 159 560
rect 225 118 255 560
rect 321 118 351 560
rect 417 118 447 560
rect 513 118 543 560
rect 609 118 639 560
rect 705 118 735 560
rect 801 118 831 560
rect -831 -560 -801 -118
rect -735 -560 -705 -118
rect -639 -560 -609 -118
rect -543 -560 -513 -118
rect -447 -560 -417 -118
rect -351 -560 -321 -118
rect -255 -560 -225 -118
rect -159 -560 -129 -118
rect -63 -560 -33 -118
rect 33 -560 63 -118
rect 129 -560 159 -118
rect 225 -560 255 -118
rect 321 -560 351 -118
rect 417 -560 447 -118
rect 513 -560 543 -118
rect 609 -560 639 -118
rect 705 -560 735 -118
rect 801 -560 831 -118
<< pdiff >>
rect -893 548 -831 560
rect -893 130 -881 548
rect -847 130 -831 548
rect -893 118 -831 130
rect -801 548 -735 560
rect -801 130 -785 548
rect -751 130 -735 548
rect -801 118 -735 130
rect -705 548 -639 560
rect -705 130 -689 548
rect -655 130 -639 548
rect -705 118 -639 130
rect -609 548 -543 560
rect -609 130 -593 548
rect -559 130 -543 548
rect -609 118 -543 130
rect -513 548 -447 560
rect -513 130 -497 548
rect -463 130 -447 548
rect -513 118 -447 130
rect -417 548 -351 560
rect -417 130 -401 548
rect -367 130 -351 548
rect -417 118 -351 130
rect -321 548 -255 560
rect -321 130 -305 548
rect -271 130 -255 548
rect -321 118 -255 130
rect -225 548 -159 560
rect -225 130 -209 548
rect -175 130 -159 548
rect -225 118 -159 130
rect -129 548 -63 560
rect -129 130 -113 548
rect -79 130 -63 548
rect -129 118 -63 130
rect -33 548 33 560
rect -33 130 -17 548
rect 17 130 33 548
rect -33 118 33 130
rect 63 548 129 560
rect 63 130 79 548
rect 113 130 129 548
rect 63 118 129 130
rect 159 548 225 560
rect 159 130 175 548
rect 209 130 225 548
rect 159 118 225 130
rect 255 548 321 560
rect 255 130 271 548
rect 305 130 321 548
rect 255 118 321 130
rect 351 548 417 560
rect 351 130 367 548
rect 401 130 417 548
rect 351 118 417 130
rect 447 548 513 560
rect 447 130 463 548
rect 497 130 513 548
rect 447 118 513 130
rect 543 548 609 560
rect 543 130 559 548
rect 593 130 609 548
rect 543 118 609 130
rect 639 548 705 560
rect 639 130 655 548
rect 689 130 705 548
rect 639 118 705 130
rect 735 548 801 560
rect 735 130 751 548
rect 785 130 801 548
rect 735 118 801 130
rect 831 548 893 560
rect 831 130 847 548
rect 881 130 893 548
rect 831 118 893 130
rect -893 -130 -831 -118
rect -893 -548 -881 -130
rect -847 -548 -831 -130
rect -893 -560 -831 -548
rect -801 -130 -735 -118
rect -801 -548 -785 -130
rect -751 -548 -735 -130
rect -801 -560 -735 -548
rect -705 -130 -639 -118
rect -705 -548 -689 -130
rect -655 -548 -639 -130
rect -705 -560 -639 -548
rect -609 -130 -543 -118
rect -609 -548 -593 -130
rect -559 -548 -543 -130
rect -609 -560 -543 -548
rect -513 -130 -447 -118
rect -513 -548 -497 -130
rect -463 -548 -447 -130
rect -513 -560 -447 -548
rect -417 -130 -351 -118
rect -417 -548 -401 -130
rect -367 -548 -351 -130
rect -417 -560 -351 -548
rect -321 -130 -255 -118
rect -321 -548 -305 -130
rect -271 -548 -255 -130
rect -321 -560 -255 -548
rect -225 -130 -159 -118
rect -225 -548 -209 -130
rect -175 -548 -159 -130
rect -225 -560 -159 -548
rect -129 -130 -63 -118
rect -129 -548 -113 -130
rect -79 -548 -63 -130
rect -129 -560 -63 -548
rect -33 -130 33 -118
rect -33 -548 -17 -130
rect 17 -548 33 -130
rect -33 -560 33 -548
rect 63 -130 129 -118
rect 63 -548 79 -130
rect 113 -548 129 -130
rect 63 -560 129 -548
rect 159 -130 225 -118
rect 159 -548 175 -130
rect 209 -548 225 -130
rect 159 -560 225 -548
rect 255 -130 321 -118
rect 255 -548 271 -130
rect 305 -548 321 -130
rect 255 -560 321 -548
rect 351 -130 417 -118
rect 351 -548 367 -130
rect 401 -548 417 -130
rect 351 -560 417 -548
rect 447 -130 513 -118
rect 447 -548 463 -130
rect 497 -548 513 -130
rect 447 -560 513 -548
rect 543 -130 609 -118
rect 543 -548 559 -130
rect 593 -548 609 -130
rect 543 -560 609 -548
rect 639 -130 705 -118
rect 639 -548 655 -130
rect 689 -548 705 -130
rect 639 -560 705 -548
rect 735 -130 801 -118
rect 735 -548 751 -130
rect 785 -548 801 -130
rect 735 -560 801 -548
rect 831 -130 893 -118
rect 831 -548 847 -130
rect 881 -548 893 -130
rect 831 -560 893 -548
<< pdiffc >>
rect -881 130 -847 548
rect -785 130 -751 548
rect -689 130 -655 548
rect -593 130 -559 548
rect -497 130 -463 548
rect -401 130 -367 548
rect -305 130 -271 548
rect -209 130 -175 548
rect -113 130 -79 548
rect -17 130 17 548
rect 79 130 113 548
rect 175 130 209 548
rect 271 130 305 548
rect 367 130 401 548
rect 463 130 497 548
rect 559 130 593 548
rect 655 130 689 548
rect 751 130 785 548
rect 847 130 881 548
rect -881 -548 -847 -130
rect -785 -548 -751 -130
rect -689 -548 -655 -130
rect -593 -548 -559 -130
rect -497 -548 -463 -130
rect -401 -548 -367 -130
rect -305 -548 -271 -130
rect -209 -548 -175 -130
rect -113 -548 -79 -130
rect -17 -548 17 -130
rect 79 -548 113 -130
rect 175 -548 209 -130
rect 271 -548 305 -130
rect 367 -548 401 -130
rect 463 -548 497 -130
rect 559 -548 593 -130
rect 655 -548 689 -130
rect 751 -548 785 -130
rect 847 -548 881 -130
<< nsubdiff >>
rect -995 709 -899 743
rect 899 709 995 743
rect -995 647 -961 709
rect 961 647 995 709
rect -995 -709 -961 -647
rect 961 -709 995 -647
rect -995 -743 -899 -709
rect 899 -743 995 -709
<< nsubdiffcont >>
rect -899 709 899 743
rect -995 -647 -961 647
rect 961 -647 995 647
rect -899 -743 899 -709
<< poly >>
rect -849 641 -783 657
rect -849 607 -833 641
rect -799 607 -783 641
rect -849 591 -783 607
rect -657 641 -591 657
rect -657 607 -641 641
rect -607 607 -591 641
rect -657 591 -591 607
rect -465 641 -399 657
rect -465 607 -449 641
rect -415 607 -399 641
rect -465 591 -399 607
rect -273 641 -207 657
rect -273 607 -257 641
rect -223 607 -207 641
rect -273 591 -207 607
rect -81 641 -15 657
rect -81 607 -65 641
rect -31 607 -15 641
rect -81 591 -15 607
rect 111 641 177 657
rect 111 607 127 641
rect 161 607 177 641
rect 111 591 177 607
rect 303 641 369 657
rect 303 607 319 641
rect 353 607 369 641
rect 303 591 369 607
rect 495 641 561 657
rect 495 607 511 641
rect 545 607 561 641
rect 495 591 561 607
rect 687 641 753 657
rect 687 607 703 641
rect 737 607 753 641
rect 687 591 753 607
rect -831 560 -801 591
rect -735 560 -705 586
rect -639 560 -609 591
rect -543 560 -513 586
rect -447 560 -417 591
rect -351 560 -321 586
rect -255 560 -225 591
rect -159 560 -129 586
rect -63 560 -33 591
rect 33 560 63 586
rect 129 560 159 591
rect 225 560 255 586
rect 321 560 351 591
rect 417 560 447 586
rect 513 560 543 591
rect 609 560 639 586
rect 705 560 735 591
rect 801 560 831 586
rect -831 92 -801 118
rect -735 87 -705 118
rect -639 92 -609 118
rect -543 87 -513 118
rect -447 92 -417 118
rect -351 87 -321 118
rect -255 92 -225 118
rect -159 87 -129 118
rect -63 92 -33 118
rect 33 87 63 118
rect 129 92 159 118
rect 225 87 255 118
rect 321 92 351 118
rect 417 87 447 118
rect 513 92 543 118
rect 609 87 639 118
rect 705 92 735 118
rect 801 87 831 118
rect -753 71 -687 87
rect -753 37 -737 71
rect -703 37 -687 71
rect -753 21 -687 37
rect -561 71 -495 87
rect -561 37 -545 71
rect -511 37 -495 71
rect -561 21 -495 37
rect -369 71 -303 87
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect 591 71 657 87
rect 591 37 607 71
rect 641 37 657 71
rect 591 21 657 37
rect 783 71 849 87
rect 783 37 799 71
rect 833 37 849 71
rect 783 21 849 37
rect -753 -37 -687 -21
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -753 -87 -687 -71
rect -561 -37 -495 -21
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -561 -87 -495 -71
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 399 -87 465 -71
rect 591 -37 657 -21
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 591 -87 657 -71
rect 783 -37 849 -21
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 783 -87 849 -71
rect -831 -118 -801 -92
rect -735 -118 -705 -87
rect -639 -118 -609 -92
rect -543 -118 -513 -87
rect -447 -118 -417 -92
rect -351 -118 -321 -87
rect -255 -118 -225 -92
rect -159 -118 -129 -87
rect -63 -118 -33 -92
rect 33 -118 63 -87
rect 129 -118 159 -92
rect 225 -118 255 -87
rect 321 -118 351 -92
rect 417 -118 447 -87
rect 513 -118 543 -92
rect 609 -118 639 -87
rect 705 -118 735 -92
rect 801 -118 831 -87
rect -831 -591 -801 -560
rect -735 -586 -705 -560
rect -639 -591 -609 -560
rect -543 -586 -513 -560
rect -447 -591 -417 -560
rect -351 -586 -321 -560
rect -255 -591 -225 -560
rect -159 -586 -129 -560
rect -63 -591 -33 -560
rect 33 -586 63 -560
rect 129 -591 159 -560
rect 225 -586 255 -560
rect 321 -591 351 -560
rect 417 -586 447 -560
rect 513 -591 543 -560
rect 609 -586 639 -560
rect 705 -591 735 -560
rect 801 -586 831 -560
rect -849 -607 -783 -591
rect -849 -641 -833 -607
rect -799 -641 -783 -607
rect -849 -657 -783 -641
rect -657 -607 -591 -591
rect -657 -641 -641 -607
rect -607 -641 -591 -607
rect -657 -657 -591 -641
rect -465 -607 -399 -591
rect -465 -641 -449 -607
rect -415 -641 -399 -607
rect -465 -657 -399 -641
rect -273 -607 -207 -591
rect -273 -641 -257 -607
rect -223 -641 -207 -607
rect -273 -657 -207 -641
rect -81 -607 -15 -591
rect -81 -641 -65 -607
rect -31 -641 -15 -607
rect -81 -657 -15 -641
rect 111 -607 177 -591
rect 111 -641 127 -607
rect 161 -641 177 -607
rect 111 -657 177 -641
rect 303 -607 369 -591
rect 303 -641 319 -607
rect 353 -641 369 -607
rect 303 -657 369 -641
rect 495 -607 561 -591
rect 495 -641 511 -607
rect 545 -641 561 -607
rect 495 -657 561 -641
rect 687 -607 753 -591
rect 687 -641 703 -607
rect 737 -641 753 -607
rect 687 -657 753 -641
<< polycont >>
rect -833 607 -799 641
rect -641 607 -607 641
rect -449 607 -415 641
rect -257 607 -223 641
rect -65 607 -31 641
rect 127 607 161 641
rect 319 607 353 641
rect 511 607 545 641
rect 703 607 737 641
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect -833 -641 -799 -607
rect -641 -641 -607 -607
rect -449 -641 -415 -607
rect -257 -641 -223 -607
rect -65 -641 -31 -607
rect 127 -641 161 -607
rect 319 -641 353 -607
rect 511 -641 545 -607
rect 703 -641 737 -607
<< locali >>
rect -995 709 -899 743
rect 899 709 995 743
rect -995 647 -961 709
rect 961 647 995 709
rect -849 607 -833 641
rect -799 607 -783 641
rect -657 607 -641 641
rect -607 607 -591 641
rect -465 607 -449 641
rect -415 607 -399 641
rect -273 607 -257 641
rect -223 607 -207 641
rect -81 607 -65 641
rect -31 607 -15 641
rect 111 607 127 641
rect 161 607 177 641
rect 303 607 319 641
rect 353 607 369 641
rect 495 607 511 641
rect 545 607 561 641
rect 687 607 703 641
rect 737 607 753 641
rect -881 548 -847 564
rect -881 114 -847 130
rect -785 548 -751 564
rect -785 114 -751 130
rect -689 548 -655 564
rect -689 114 -655 130
rect -593 548 -559 564
rect -593 114 -559 130
rect -497 548 -463 564
rect -497 114 -463 130
rect -401 548 -367 564
rect -401 114 -367 130
rect -305 548 -271 564
rect -305 114 -271 130
rect -209 548 -175 564
rect -209 114 -175 130
rect -113 548 -79 564
rect -113 114 -79 130
rect -17 548 17 564
rect -17 114 17 130
rect 79 548 113 564
rect 79 114 113 130
rect 175 548 209 564
rect 175 114 209 130
rect 271 548 305 564
rect 271 114 305 130
rect 367 548 401 564
rect 367 114 401 130
rect 463 548 497 564
rect 463 114 497 130
rect 559 548 593 564
rect 559 114 593 130
rect 655 548 689 564
rect 655 114 689 130
rect 751 548 785 564
rect 751 114 785 130
rect 847 548 881 564
rect 847 114 881 130
rect -753 37 -737 71
rect -703 37 -687 71
rect -561 37 -545 71
rect -511 37 -495 71
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect 591 37 607 71
rect 641 37 657 71
rect 783 37 799 71
rect 833 37 849 71
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 783 -71 799 -37
rect 833 -71 849 -37
rect -881 -130 -847 -114
rect -881 -564 -847 -548
rect -785 -130 -751 -114
rect -785 -564 -751 -548
rect -689 -130 -655 -114
rect -689 -564 -655 -548
rect -593 -130 -559 -114
rect -593 -564 -559 -548
rect -497 -130 -463 -114
rect -497 -564 -463 -548
rect -401 -130 -367 -114
rect -401 -564 -367 -548
rect -305 -130 -271 -114
rect -305 -564 -271 -548
rect -209 -130 -175 -114
rect -209 -564 -175 -548
rect -113 -130 -79 -114
rect -113 -564 -79 -548
rect -17 -130 17 -114
rect -17 -564 17 -548
rect 79 -130 113 -114
rect 79 -564 113 -548
rect 175 -130 209 -114
rect 175 -564 209 -548
rect 271 -130 305 -114
rect 271 -564 305 -548
rect 367 -130 401 -114
rect 367 -564 401 -548
rect 463 -130 497 -114
rect 463 -564 497 -548
rect 559 -130 593 -114
rect 559 -564 593 -548
rect 655 -130 689 -114
rect 655 -564 689 -548
rect 751 -130 785 -114
rect 751 -564 785 -548
rect 847 -130 881 -114
rect 847 -564 881 -548
rect -849 -641 -833 -607
rect -799 -641 -783 -607
rect -657 -641 -641 -607
rect -607 -641 -591 -607
rect -465 -641 -449 -607
rect -415 -641 -399 -607
rect -273 -641 -257 -607
rect -223 -641 -207 -607
rect -81 -641 -65 -607
rect -31 -641 -15 -607
rect 111 -641 127 -607
rect 161 -641 177 -607
rect 303 -641 319 -607
rect 353 -641 369 -607
rect 495 -641 511 -607
rect 545 -641 561 -607
rect 687 -641 703 -607
rect 737 -641 753 -607
rect -995 -709 -961 -647
rect 961 -709 995 -647
rect -995 -743 -899 -709
rect 899 -743 995 -709
<< viali >>
rect -833 607 -799 641
rect -641 607 -607 641
rect -449 607 -415 641
rect -257 607 -223 641
rect -65 607 -31 641
rect 127 607 161 641
rect 319 607 353 641
rect 511 607 545 641
rect 703 607 737 641
rect -881 130 -847 548
rect -785 130 -751 548
rect -689 130 -655 548
rect -593 130 -559 548
rect -497 130 -463 548
rect -401 130 -367 548
rect -305 130 -271 548
rect -209 130 -175 548
rect -113 130 -79 548
rect -17 130 17 548
rect 79 130 113 548
rect 175 130 209 548
rect 271 130 305 548
rect 367 130 401 548
rect 463 130 497 548
rect 559 130 593 548
rect 655 130 689 548
rect 751 130 785 548
rect 847 130 881 548
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect -881 -548 -847 -130
rect -785 -548 -751 -130
rect -689 -548 -655 -130
rect -593 -548 -559 -130
rect -497 -548 -463 -130
rect -401 -548 -367 -130
rect -305 -548 -271 -130
rect -209 -548 -175 -130
rect -113 -548 -79 -130
rect -17 -548 17 -130
rect 79 -548 113 -130
rect 175 -548 209 -130
rect 271 -548 305 -130
rect 367 -548 401 -130
rect 463 -548 497 -130
rect 559 -548 593 -130
rect 655 -548 689 -130
rect 751 -548 785 -130
rect 847 -548 881 -130
rect -833 -641 -799 -607
rect -641 -641 -607 -607
rect -449 -641 -415 -607
rect -257 -641 -223 -607
rect -65 -641 -31 -607
rect 127 -641 161 -607
rect 319 -641 353 -607
rect 511 -641 545 -607
rect 703 -641 737 -607
<< metal1 >>
rect -845 641 -787 647
rect -845 607 -833 641
rect -799 607 -787 641
rect -845 601 -787 607
rect -653 641 -595 647
rect -653 607 -641 641
rect -607 607 -595 641
rect -653 601 -595 607
rect -461 641 -403 647
rect -461 607 -449 641
rect -415 607 -403 641
rect -461 601 -403 607
rect -269 641 -211 647
rect -269 607 -257 641
rect -223 607 -211 641
rect -269 601 -211 607
rect -77 641 -19 647
rect -77 607 -65 641
rect -31 607 -19 641
rect -77 601 -19 607
rect 115 641 173 647
rect 115 607 127 641
rect 161 607 173 641
rect 115 601 173 607
rect 307 641 365 647
rect 307 607 319 641
rect 353 607 365 641
rect 307 601 365 607
rect 499 641 557 647
rect 499 607 511 641
rect 545 607 557 641
rect 499 601 557 607
rect 691 641 749 647
rect 691 607 703 641
rect 737 607 749 641
rect 691 601 749 607
rect -887 548 -841 560
rect -887 130 -881 548
rect -847 130 -841 548
rect -887 118 -841 130
rect -791 548 -745 560
rect -791 130 -785 548
rect -751 130 -745 548
rect -791 118 -745 130
rect -695 548 -649 560
rect -695 130 -689 548
rect -655 130 -649 548
rect -695 118 -649 130
rect -599 548 -553 560
rect -599 130 -593 548
rect -559 130 -553 548
rect -599 118 -553 130
rect -503 548 -457 560
rect -503 130 -497 548
rect -463 130 -457 548
rect -503 118 -457 130
rect -407 548 -361 560
rect -407 130 -401 548
rect -367 130 -361 548
rect -407 118 -361 130
rect -311 548 -265 560
rect -311 130 -305 548
rect -271 130 -265 548
rect -311 118 -265 130
rect -215 548 -169 560
rect -215 130 -209 548
rect -175 130 -169 548
rect -215 118 -169 130
rect -119 548 -73 560
rect -119 130 -113 548
rect -79 130 -73 548
rect -119 118 -73 130
rect -23 548 23 560
rect -23 130 -17 548
rect 17 130 23 548
rect -23 118 23 130
rect 73 548 119 560
rect 73 130 79 548
rect 113 130 119 548
rect 73 118 119 130
rect 169 548 215 560
rect 169 130 175 548
rect 209 130 215 548
rect 169 118 215 130
rect 265 548 311 560
rect 265 130 271 548
rect 305 130 311 548
rect 265 118 311 130
rect 361 548 407 560
rect 361 130 367 548
rect 401 130 407 548
rect 361 118 407 130
rect 457 548 503 560
rect 457 130 463 548
rect 497 130 503 548
rect 457 118 503 130
rect 553 548 599 560
rect 553 130 559 548
rect 593 130 599 548
rect 553 118 599 130
rect 649 548 695 560
rect 649 130 655 548
rect 689 130 695 548
rect 649 118 695 130
rect 745 548 791 560
rect 745 130 751 548
rect 785 130 791 548
rect 745 118 791 130
rect 841 548 887 560
rect 841 130 847 548
rect 881 130 887 548
rect 841 118 887 130
rect -749 71 -691 77
rect -749 37 -737 71
rect -703 37 -691 71
rect -749 31 -691 37
rect -557 71 -499 77
rect -557 37 -545 71
rect -511 37 -499 71
rect -557 31 -499 37
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect 595 71 653 77
rect 595 37 607 71
rect 641 37 653 71
rect 595 31 653 37
rect 787 71 845 77
rect 787 37 799 71
rect 833 37 845 71
rect 787 31 845 37
rect -749 -37 -691 -31
rect -749 -71 -737 -37
rect -703 -71 -691 -37
rect -749 -77 -691 -71
rect -557 -37 -499 -31
rect -557 -71 -545 -37
rect -511 -71 -499 -37
rect -557 -77 -499 -71
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect 595 -37 653 -31
rect 595 -71 607 -37
rect 641 -71 653 -37
rect 595 -77 653 -71
rect 787 -37 845 -31
rect 787 -71 799 -37
rect 833 -71 845 -37
rect 787 -77 845 -71
rect -887 -130 -841 -118
rect -887 -548 -881 -130
rect -847 -548 -841 -130
rect -887 -560 -841 -548
rect -791 -130 -745 -118
rect -791 -548 -785 -130
rect -751 -548 -745 -130
rect -791 -560 -745 -548
rect -695 -130 -649 -118
rect -695 -548 -689 -130
rect -655 -548 -649 -130
rect -695 -560 -649 -548
rect -599 -130 -553 -118
rect -599 -548 -593 -130
rect -559 -548 -553 -130
rect -599 -560 -553 -548
rect -503 -130 -457 -118
rect -503 -548 -497 -130
rect -463 -548 -457 -130
rect -503 -560 -457 -548
rect -407 -130 -361 -118
rect -407 -548 -401 -130
rect -367 -548 -361 -130
rect -407 -560 -361 -548
rect -311 -130 -265 -118
rect -311 -548 -305 -130
rect -271 -548 -265 -130
rect -311 -560 -265 -548
rect -215 -130 -169 -118
rect -215 -548 -209 -130
rect -175 -548 -169 -130
rect -215 -560 -169 -548
rect -119 -130 -73 -118
rect -119 -548 -113 -130
rect -79 -548 -73 -130
rect -119 -560 -73 -548
rect -23 -130 23 -118
rect -23 -548 -17 -130
rect 17 -548 23 -130
rect -23 -560 23 -548
rect 73 -130 119 -118
rect 73 -548 79 -130
rect 113 -548 119 -130
rect 73 -560 119 -548
rect 169 -130 215 -118
rect 169 -548 175 -130
rect 209 -548 215 -130
rect 169 -560 215 -548
rect 265 -130 311 -118
rect 265 -548 271 -130
rect 305 -548 311 -130
rect 265 -560 311 -548
rect 361 -130 407 -118
rect 361 -548 367 -130
rect 401 -548 407 -130
rect 361 -560 407 -548
rect 457 -130 503 -118
rect 457 -548 463 -130
rect 497 -548 503 -130
rect 457 -560 503 -548
rect 553 -130 599 -118
rect 553 -548 559 -130
rect 593 -548 599 -130
rect 553 -560 599 -548
rect 649 -130 695 -118
rect 649 -548 655 -130
rect 689 -548 695 -130
rect 649 -560 695 -548
rect 745 -130 791 -118
rect 745 -548 751 -130
rect 785 -548 791 -130
rect 745 -560 791 -548
rect 841 -130 887 -118
rect 841 -548 847 -130
rect 881 -548 887 -130
rect 841 -560 887 -548
rect -845 -607 -787 -601
rect -845 -641 -833 -607
rect -799 -641 -787 -607
rect -845 -647 -787 -641
rect -653 -607 -595 -601
rect -653 -641 -641 -607
rect -607 -641 -595 -607
rect -653 -647 -595 -641
rect -461 -607 -403 -601
rect -461 -641 -449 -607
rect -415 -641 -403 -607
rect -461 -647 -403 -641
rect -269 -607 -211 -601
rect -269 -641 -257 -607
rect -223 -641 -211 -607
rect -269 -647 -211 -641
rect -77 -607 -19 -601
rect -77 -641 -65 -607
rect -31 -641 -19 -607
rect -77 -647 -19 -641
rect 115 -607 173 -601
rect 115 -641 127 -607
rect 161 -641 173 -607
rect 115 -647 173 -641
rect 307 -607 365 -601
rect 307 -641 319 -607
rect 353 -641 365 -607
rect 307 -647 365 -641
rect 499 -607 557 -601
rect 499 -641 511 -607
rect 545 -641 557 -607
rect 499 -647 557 -641
rect 691 -607 749 -601
rect 691 -641 703 -607
rect 737 -641 749 -607
rect 691 -647 749 -641
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -978 -726 978 726
string parameters w 2.21 l 0.15 m 2 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
