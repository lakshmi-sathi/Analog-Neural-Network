magic
tech sky130A
magscale 1 2
timestamp 1627111729
<< xpolycontact >>
rect -141 59 141 491
rect -141 -491 141 -59
<< xpolyres >>
rect -141 -59 141 59
<< viali >>
rect -125 76 125 473
rect -125 -473 125 -76
<< metal1 >>
rect -131 473 131 485
rect -131 76 -125 473
rect 125 76 131 473
rect -131 64 131 76
rect -131 -76 131 -64
rect -131 -473 -125 -76
rect 125 -473 131 -76
rect -131 -485 131 -473
<< res1p41 >>
rect -143 -61 143 61
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string parameters w 1.410 l 0.59 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 1.007k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
