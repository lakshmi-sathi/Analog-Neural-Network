magic
tech sky130A
magscale 1 2
timestamp 1627921586
<< xpolycontact >>
rect -35 292 35 724
rect -35 -724 35 -292
<< ppolyres >>
rect -35 -292 35 292
<< viali >>
rect -19 309 19 706
rect -19 -706 19 -309
<< metal1 >>
rect -25 706 25 718
rect -25 309 -19 706
rect 19 309 25 706
rect -25 297 25 309
rect -25 -309 25 -297
rect -25 -706 -19 -309
rect 19 -706 25 -309
rect -25 -718 25 -706
<< res0p35 >>
rect -37 -294 37 294
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string parameters w 0.350 l 2.92 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 2.777k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 0.350 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
