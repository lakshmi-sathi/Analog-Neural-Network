magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 76 35 508
rect -35 -508 35 -76
<< xpolyres >>
rect -35 -76 35 76
<< viali >>
rect -17 454 17 488
rect -17 382 17 416
rect -17 310 17 344
rect -17 238 17 272
rect -17 166 17 200
rect -17 94 17 128
rect -17 -129 17 -95
rect -17 -201 17 -167
rect -17 -273 17 -239
rect -17 -345 17 -311
rect -17 -417 17 -383
rect -17 -489 17 -455
<< metal1 >>
rect -25 488 25 502
rect -25 454 -17 488
rect 17 454 25 488
rect -25 416 25 454
rect -25 382 -17 416
rect 17 382 25 416
rect -25 344 25 382
rect -25 310 -17 344
rect 17 310 25 344
rect -25 272 25 310
rect -25 238 -17 272
rect 17 238 25 272
rect -25 200 25 238
rect -25 166 -17 200
rect 17 166 25 200
rect -25 128 25 166
rect -25 94 -17 128
rect 17 94 25 128
rect -25 81 25 94
rect -25 -95 25 -81
rect -25 -129 -17 -95
rect 17 -129 25 -95
rect -25 -167 25 -129
rect -25 -201 -17 -167
rect 17 -201 25 -167
rect -25 -239 25 -201
rect -25 -273 -17 -239
rect 17 -273 25 -239
rect -25 -311 25 -273
rect -25 -345 -17 -311
rect 17 -345 25 -311
rect -25 -383 25 -345
rect -25 -417 -17 -383
rect 17 -417 25 -383
rect -25 -455 25 -417
rect -25 -489 -17 -455
rect 17 -489 25 -455
rect -25 -502 25 -489
<< end >>
