magic
tech sky130A
magscale 1 2
timestamp 1628066849
<< error_p >>
rect -29 959 29 965
rect -29 925 -17 959
rect -29 919 29 925
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
<< pwell >>
rect -211 -1097 211 1097
<< nmos >>
rect -15 47 15 887
rect -15 -949 15 -109
<< ndiff >>
rect -73 875 -15 887
rect -73 59 -61 875
rect -27 59 -15 875
rect -73 47 -15 59
rect 15 875 73 887
rect 15 59 27 875
rect 61 59 73 875
rect 15 47 73 59
rect -73 -121 -15 -109
rect -73 -937 -61 -121
rect -27 -937 -15 -121
rect -73 -949 -15 -937
rect 15 -121 73 -109
rect 15 -937 27 -121
rect 61 -937 73 -121
rect 15 -949 73 -937
<< ndiffc >>
rect -61 59 -27 875
rect 27 59 61 875
rect -61 -937 -27 -121
rect 27 -937 61 -121
<< psubdiff >>
rect -175 1027 -79 1061
rect 79 1027 175 1061
rect -175 965 -141 1027
rect 141 965 175 1027
rect -175 -1027 -141 -965
rect 141 -1027 175 -965
rect -175 -1061 -79 -1027
rect 79 -1061 175 -1027
<< psubdiffcont >>
rect -79 1027 79 1061
rect -175 -965 -141 965
rect 141 -965 175 965
rect -79 -1061 79 -1027
<< poly >>
rect -33 959 33 975
rect -33 925 -17 959
rect 17 925 33 959
rect -33 909 33 925
rect -15 887 15 909
rect -15 21 15 47
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -975 15 -949
<< polycont >>
rect -17 925 17 959
rect -17 -71 17 -37
<< locali >>
rect -175 1027 -79 1061
rect 79 1027 175 1061
rect -175 965 -141 1027
rect 141 965 175 1027
rect -33 925 -17 959
rect 17 925 33 959
rect -61 875 -27 891
rect -61 43 -27 59
rect 27 875 61 891
rect 27 43 61 59
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -953 -27 -937
rect 27 -121 61 -105
rect 27 -953 61 -937
rect -175 -1027 -141 -965
rect 141 -1027 175 -965
rect -175 -1061 -79 -1027
rect 79 -1061 175 -1027
<< viali >>
rect -17 925 17 959
rect -61 59 -27 875
rect 27 59 61 875
rect -17 -71 17 -37
rect -61 -937 -27 -121
rect 27 -937 61 -121
<< metal1 >>
rect -29 959 29 965
rect -29 925 -17 959
rect 17 925 29 959
rect -29 919 29 925
rect -67 875 -21 887
rect -67 59 -61 875
rect -27 59 -21 875
rect -67 47 -21 59
rect 21 875 67 887
rect 21 59 27 875
rect 61 59 67 875
rect 21 47 67 59
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -937 -61 -121
rect -27 -937 -21 -121
rect -67 -949 -21 -937
rect 21 -121 67 -109
rect 21 -937 27 -121
rect 61 -937 67 -121
rect 21 -949 67 -937
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -1044 158 1044
string parameters w 4.2 l 0.150 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
