magic
tech sky130A
magscale 1 2
timestamp 1627923075
<< xpolycontact >>
rect -35 280 35 712
rect -35 -712 35 -280
<< xpolyres >>
rect -35 -280 35 280
<< viali >>
rect -19 297 19 694
rect -19 -694 19 -297
<< metal1 >>
rect -25 694 25 706
rect -25 297 -19 694
rect 19 297 25 694
rect -25 285 25 297
rect -25 -297 25 -285
rect -25 -694 -19 -297
rect 19 -694 25 -297
rect -25 -706 25 -694
<< res0p35 >>
rect -37 -282 37 282
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 2.8 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 16.685k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
