magic
tech sky130A
magscale 1 2
timestamp 1627805142
<< xpolycontact >>
rect -35 75 35 507
rect -35 -507 35 -75
<< xpolyres >>
rect -35 -75 35 75
<< viali >>
rect -19 92 19 489
rect -19 -489 19 -92
<< metal1 >>
rect -25 489 25 501
rect -25 92 -19 489
rect 19 92 25 489
rect -25 80 25 92
rect -25 -92 25 -80
rect -25 -489 -19 -92
rect 19 -489 25 -92
rect -25 -501 25 -489
<< res0p35 >>
rect -37 -77 37 77
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 0.75 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 4.971k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
