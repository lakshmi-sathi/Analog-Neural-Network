magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< locali >>
rect 126 1627 224 1630
rect 126 1593 158 1627
rect 192 1593 224 1627
rect 126 1555 224 1593
rect 126 1521 158 1555
rect 192 1521 224 1555
rect 126 1483 224 1521
rect 126 1449 158 1483
rect 192 1449 224 1483
rect 126 1411 224 1449
rect 126 1377 158 1411
rect 192 1377 224 1411
rect 126 1339 224 1377
rect 126 1305 158 1339
rect 192 1305 224 1339
rect 126 1267 224 1305
rect 126 1233 158 1267
rect 192 1233 224 1267
rect 126 1195 224 1233
rect 126 1161 158 1195
rect 192 1161 224 1195
rect 126 1123 224 1161
rect 2558 1138 2565 1160
rect 126 1089 158 1123
rect 192 1089 224 1123
rect 126 1051 224 1089
rect 126 1017 158 1051
rect 192 1017 224 1051
rect 126 979 224 1017
rect 2479 1125 2513 1129
rect 2527 1125 2561 1131
rect 2479 1012 2561 1125
rect 126 945 158 979
rect 192 945 224 979
rect 2190 978 2561 1012
rect 126 907 224 945
rect 126 873 158 907
rect 192 873 224 907
rect 126 835 224 873
rect 126 801 158 835
rect 192 801 224 835
rect 126 763 224 801
rect 126 729 158 763
rect 192 729 224 763
rect 126 726 224 729
rect 8149 200 8369 234
rect 8165 173 8369 200
rect 8335 102 8369 173
rect 8334 18 8530 102
<< viali >>
rect 158 1593 192 1627
rect 158 1521 192 1555
rect 158 1449 192 1483
rect 158 1377 192 1411
rect 158 1305 192 1339
rect 158 1233 192 1267
rect 158 1161 192 1195
rect 158 1089 192 1123
rect 158 1017 192 1051
rect 158 945 192 979
rect 158 873 192 907
rect 158 801 192 835
rect 158 729 192 763
<< metal1 >>
rect 2316 2400 2960 2430
rect 2316 2374 3294 2400
rect 134 1650 236 1654
rect 108 1632 236 1650
rect 108 1627 270 1632
rect 108 1593 158 1627
rect 192 1593 270 1627
rect 108 1555 270 1593
rect 108 1521 158 1555
rect 192 1521 270 1555
rect 108 1483 270 1521
rect 108 1449 158 1483
rect 192 1449 270 1483
rect 2316 1450 2456 2374
rect 2816 2352 3294 2374
rect 2816 2350 2958 2352
rect 108 1411 270 1449
rect 108 1377 158 1411
rect 192 1377 270 1411
rect 108 1339 270 1377
rect 108 1305 158 1339
rect 192 1305 270 1339
rect 108 1267 270 1305
rect 108 1233 158 1267
rect 192 1233 270 1267
rect 108 1195 270 1233
rect 108 1161 158 1195
rect 192 1161 270 1195
rect 108 1123 270 1161
rect 108 1108 158 1123
rect -762 1089 158 1108
rect 192 1108 270 1123
rect 2250 1404 2456 1450
rect 2250 1352 2303 1404
rect 2355 1352 2456 1404
rect 2250 1340 2456 1352
rect 2250 1288 2303 1340
rect 2355 1288 2456 1340
rect 2250 1276 2456 1288
rect 2250 1224 2303 1276
rect 2355 1270 2456 1276
rect 3956 1378 4044 1384
rect 4246 1378 4300 1992
rect 4429 1378 4483 1989
rect 4623 1378 4677 1981
rect 4823 1378 4877 1969
rect 5011 1378 5065 1969
rect 5207 1378 5261 1963
rect 5387 1378 5441 1985
rect 5583 1378 5637 1963
rect 5779 1378 5833 1965
rect 5975 1378 6029 1967
rect 6155 1378 6209 1969
rect 6355 1378 6409 1969
rect 6551 1378 6605 1977
rect 6739 1378 6793 1973
rect 7754 1491 7948 1492
rect 8260 1491 8443 1493
rect 7754 1474 8443 1491
rect 7390 1453 8443 1474
rect 7390 1426 7948 1453
rect 3956 1368 6834 1378
rect 2355 1224 2498 1270
rect 3956 1252 3994 1368
rect 6798 1252 6834 1368
rect 3956 1242 6834 1252
rect 3956 1236 4094 1242
rect 2250 1212 2498 1224
rect 2250 1160 2303 1212
rect 2355 1182 2498 1212
rect 2355 1160 2412 1182
rect 2250 1114 2412 1160
rect 192 1089 352 1108
rect -762 1051 352 1089
rect -762 1017 158 1051
rect 192 1017 352 1051
rect -762 979 352 1017
rect -762 945 158 979
rect 192 945 352 979
rect -762 907 352 945
rect -762 873 158 907
rect 192 873 352 907
rect -762 835 352 873
rect -762 801 158 835
rect 192 801 352 835
rect -1354 382 -932 776
rect -762 763 352 801
rect -762 729 158 763
rect 192 729 352 763
rect 4042 744 4094 1236
rect 4234 744 4286 1242
rect 4430 744 4482 1242
rect 4614 744 4666 1242
rect 4806 744 4858 1242
rect 5004 744 5056 1242
rect 5196 744 5248 1242
rect 5388 744 5440 1242
rect 5580 744 5632 1242
rect 5776 744 5828 1242
rect 5964 744 6016 1242
rect 6160 744 6212 1242
rect 6344 744 6396 1242
rect 8260 936 8443 1453
rect 8260 894 8444 936
rect -762 710 352 729
rect -306 706 210 710
rect 8260 586 8298 894
rect 8414 586 8444 894
rect 10412 686 10656 1630
rect -1346 -46 -924 118
rect -762 60 -340 454
rect 8260 400 8444 586
rect 8258 344 8444 400
rect 8224 256 8444 344
rect -10 234 166 238
rect -194 218 166 234
rect -194 -26 20 218
rect 136 -26 166 218
rect -194 -46 166 -26
rect -1346 -54 78 -46
rect -1346 -142 -32 -54
<< via1 >>
rect 2303 1352 2355 1404
rect 2303 1288 2355 1340
rect 2303 1224 2355 1276
rect 3994 1252 6798 1368
rect 2303 1160 2355 1212
rect 8298 586 8414 894
rect 20 -26 136 218
<< metal2 >>
rect 66 2780 10696 2910
rect 254 2666 2318 2780
rect 2455 2560 4030 2680
rect 2455 2559 3822 2560
rect 3880 1947 4030 2560
rect 3880 1797 4032 1947
rect 3881 1760 4032 1797
rect 4156 1760 8268 1762
rect 3881 1712 8268 1760
rect 3881 1656 4130 1712
rect 4186 1656 4210 1712
rect 4266 1656 4290 1712
rect 4346 1656 4370 1712
rect 4426 1656 4450 1712
rect 4506 1656 4530 1712
rect 4586 1656 4610 1712
rect 4666 1656 4690 1712
rect 4746 1656 4770 1712
rect 4826 1656 4850 1712
rect 4906 1656 4930 1712
rect 4986 1656 5010 1712
rect 5066 1656 5090 1712
rect 5146 1656 5170 1712
rect 5226 1656 5250 1712
rect 5306 1656 5330 1712
rect 5386 1656 5410 1712
rect 5466 1656 5490 1712
rect 5546 1656 5570 1712
rect 5626 1656 5650 1712
rect 5706 1656 5730 1712
rect 5786 1656 5810 1712
rect 5866 1656 5890 1712
rect 5946 1656 5970 1712
rect 6026 1656 6050 1712
rect 6106 1656 6130 1712
rect 6186 1656 6210 1712
rect 6266 1656 6290 1712
rect 6346 1656 6370 1712
rect 6426 1656 6450 1712
rect 6506 1656 6530 1712
rect 6586 1656 6610 1712
rect 6666 1656 6690 1712
rect 6746 1656 6770 1712
rect 6826 1656 6850 1712
rect 6906 1656 6930 1712
rect 6986 1656 7010 1712
rect 7066 1656 7090 1712
rect 7146 1656 7170 1712
rect 7226 1656 7250 1712
rect 7306 1656 7330 1712
rect 7386 1656 7410 1712
rect 7466 1656 7490 1712
rect 7546 1656 7570 1712
rect 7626 1656 7650 1712
rect 7706 1656 7730 1712
rect 7786 1656 7810 1712
rect 7866 1656 7890 1712
rect 7946 1656 7970 1712
rect 8026 1656 8050 1712
rect 8106 1656 8130 1712
rect 8186 1656 8268 1712
rect 3881 1612 8268 1656
rect 3881 1611 4143 1612
rect 3881 1609 4031 1611
rect 2258 1429 2400 1444
rect 2258 1373 2302 1429
rect 2358 1373 2400 1429
rect 2258 1352 2303 1373
rect 2355 1352 2400 1373
rect 2258 1349 2400 1352
rect 2258 1293 2302 1349
rect 2358 1293 2400 1349
rect 2258 1288 2303 1293
rect 2355 1288 2400 1293
rect 2258 1276 2400 1288
rect 2258 1269 2303 1276
rect 2355 1269 2400 1276
rect 2258 1213 2302 1269
rect 2358 1213 2400 1269
rect 3962 1378 6824 1388
rect 3962 1242 3968 1378
rect 3962 1232 6824 1242
rect 2258 1212 2400 1213
rect 2258 1189 2303 1212
rect 2355 1189 2400 1212
rect 2258 1133 2302 1189
rect 2358 1133 2400 1189
rect 2258 1120 2400 1133
rect 3708 1054 3812 1084
rect 4006 1054 6848 1064
rect 3708 1018 6848 1054
rect 3708 962 4020 1018
rect 4076 962 4100 1018
rect 4156 962 4180 1018
rect 4236 962 4260 1018
rect 4316 962 4340 1018
rect 4396 962 4420 1018
rect 4476 962 4500 1018
rect 4556 962 4580 1018
rect 4636 962 4660 1018
rect 4716 962 4740 1018
rect 4796 962 4820 1018
rect 4876 962 4900 1018
rect 4956 962 4980 1018
rect 5036 962 5060 1018
rect 5116 962 5140 1018
rect 5196 962 5220 1018
rect 5276 962 5300 1018
rect 5356 962 5380 1018
rect 5436 962 5460 1018
rect 5516 962 5540 1018
rect 5596 962 5620 1018
rect 5676 962 5700 1018
rect 5756 962 5780 1018
rect 5836 962 5860 1018
rect 5916 962 5940 1018
rect 5996 962 6020 1018
rect 6076 962 6100 1018
rect 6156 962 6180 1018
rect 6236 962 6260 1018
rect 6316 962 6340 1018
rect 6396 962 6420 1018
rect 6476 962 6500 1018
rect 6556 962 6580 1018
rect 6636 962 6848 1018
rect 3708 926 6848 962
rect 4006 918 6848 926
rect 0 218 156 248
rect 0 204 20 218
rect 136 204 156 218
rect 0 -12 10 204
rect 146 -12 156 204
rect 6701 197 6847 918
rect 8276 894 8434 906
rect 8276 586 8298 894
rect 8414 586 8434 894
rect 8276 570 8434 586
rect 6701 146 6850 197
rect 6701 141 6868 146
rect 6701 51 8240 141
rect 6702 -5 8240 51
rect 6702 -8 6888 -5
rect 0 -26 20 -12
rect 136 -26 156 -12
rect 0 -56 156 -26
rect 94 -234 10724 -104
<< via2 >>
rect 4130 1656 4186 1712
rect 4210 1656 4266 1712
rect 4290 1656 4346 1712
rect 4370 1656 4426 1712
rect 4450 1656 4506 1712
rect 4530 1656 4586 1712
rect 4610 1656 4666 1712
rect 4690 1656 4746 1712
rect 4770 1656 4826 1712
rect 4850 1656 4906 1712
rect 4930 1656 4986 1712
rect 5010 1656 5066 1712
rect 5090 1656 5146 1712
rect 5170 1656 5226 1712
rect 5250 1656 5306 1712
rect 5330 1656 5386 1712
rect 5410 1656 5466 1712
rect 5490 1656 5546 1712
rect 5570 1656 5626 1712
rect 5650 1656 5706 1712
rect 5730 1656 5786 1712
rect 5810 1656 5866 1712
rect 5890 1656 5946 1712
rect 5970 1656 6026 1712
rect 6050 1656 6106 1712
rect 6130 1656 6186 1712
rect 6210 1656 6266 1712
rect 6290 1656 6346 1712
rect 6370 1656 6426 1712
rect 6450 1656 6506 1712
rect 6530 1656 6586 1712
rect 6610 1656 6666 1712
rect 6690 1656 6746 1712
rect 6770 1656 6826 1712
rect 6850 1656 6906 1712
rect 6930 1656 6986 1712
rect 7010 1656 7066 1712
rect 7090 1656 7146 1712
rect 7170 1656 7226 1712
rect 7250 1656 7306 1712
rect 7330 1656 7386 1712
rect 7410 1656 7466 1712
rect 7490 1656 7546 1712
rect 7570 1656 7626 1712
rect 7650 1656 7706 1712
rect 7730 1656 7786 1712
rect 7810 1656 7866 1712
rect 7890 1656 7946 1712
rect 7970 1656 8026 1712
rect 8050 1656 8106 1712
rect 8130 1656 8186 1712
rect 2302 1404 2358 1429
rect 2302 1373 2303 1404
rect 2303 1373 2355 1404
rect 2355 1373 2358 1404
rect 2302 1340 2358 1349
rect 2302 1293 2303 1340
rect 2303 1293 2355 1340
rect 2355 1293 2358 1340
rect 2302 1224 2303 1269
rect 2303 1224 2355 1269
rect 2355 1224 2358 1269
rect 2302 1213 2358 1224
rect 3968 1368 6824 1378
rect 3968 1252 3994 1368
rect 3994 1252 6798 1368
rect 6798 1252 6824 1368
rect 3968 1242 6824 1252
rect 2302 1160 2303 1189
rect 2303 1160 2355 1189
rect 2355 1160 2358 1189
rect 2302 1133 2358 1160
rect 4020 962 4076 1018
rect 4100 962 4156 1018
rect 4180 962 4236 1018
rect 4260 962 4316 1018
rect 4340 962 4396 1018
rect 4420 962 4476 1018
rect 4500 962 4556 1018
rect 4580 962 4636 1018
rect 4660 962 4716 1018
rect 4740 962 4796 1018
rect 4820 962 4876 1018
rect 4900 962 4956 1018
rect 4980 962 5036 1018
rect 5060 962 5116 1018
rect 5140 962 5196 1018
rect 5220 962 5276 1018
rect 5300 962 5356 1018
rect 5380 962 5436 1018
rect 5460 962 5516 1018
rect 5540 962 5596 1018
rect 5620 962 5676 1018
rect 5700 962 5756 1018
rect 5780 962 5836 1018
rect 5860 962 5916 1018
rect 5940 962 5996 1018
rect 6020 962 6076 1018
rect 6100 962 6156 1018
rect 6180 962 6236 1018
rect 6260 962 6316 1018
rect 6340 962 6396 1018
rect 6420 962 6476 1018
rect 6500 962 6556 1018
rect 6580 962 6636 1018
rect 10 -12 20 204
rect 20 -12 136 204
rect 136 -12 146 204
rect 8325 793 8381 849
rect 8325 713 8381 769
rect 8325 633 8381 689
<< metal3 >>
rect 4162 1760 8274 1846
rect 4068 1712 8274 1760
rect 4068 1656 4130 1712
rect 4186 1656 4210 1712
rect 4266 1656 4290 1712
rect 4346 1656 4370 1712
rect 4426 1656 4450 1712
rect 4506 1656 4530 1712
rect 4586 1656 4610 1712
rect 4666 1656 4690 1712
rect 4746 1656 4770 1712
rect 4826 1656 4850 1712
rect 4906 1656 4930 1712
rect 4986 1656 5010 1712
rect 5066 1656 5090 1712
rect 5146 1656 5170 1712
rect 5226 1656 5250 1712
rect 5306 1656 5330 1712
rect 5386 1656 5410 1712
rect 5466 1656 5490 1712
rect 5546 1656 5570 1712
rect 5626 1656 5650 1712
rect 5706 1656 5730 1712
rect 5786 1656 5810 1712
rect 5866 1656 5890 1712
rect 5946 1656 5970 1712
rect 6026 1656 6050 1712
rect 6106 1656 6130 1712
rect 6186 1656 6210 1712
rect 6266 1656 6290 1712
rect 6346 1656 6370 1712
rect 6426 1656 6450 1712
rect 6506 1656 6530 1712
rect 6586 1656 6610 1712
rect 6666 1656 6690 1712
rect 6746 1656 6770 1712
rect 6826 1656 6850 1712
rect 6906 1656 6930 1712
rect 6986 1656 7010 1712
rect 7066 1656 7090 1712
rect 7146 1656 7170 1712
rect 7226 1656 7250 1712
rect 7306 1656 7330 1712
rect 7386 1656 7410 1712
rect 7466 1656 7490 1712
rect 7546 1656 7570 1712
rect 7626 1656 7650 1712
rect 7706 1656 7730 1712
rect 7786 1656 7810 1712
rect 7866 1656 7890 1712
rect 7946 1656 7970 1712
rect 8026 1656 8050 1712
rect 8106 1656 8130 1712
rect 8186 1688 8274 1712
rect 8186 1656 8264 1688
rect 4068 1608 8264 1656
rect 2182 1429 2400 1480
rect 2182 1373 2302 1429
rect 2358 1373 2400 1429
rect 2182 1349 2400 1373
rect 3902 1383 4044 1384
rect 3902 1378 6834 1383
rect 3902 1362 3968 1378
rect 2182 1293 2302 1349
rect 2358 1293 2400 1349
rect 2182 1269 2400 1293
rect 2182 1213 2302 1269
rect 2358 1213 2400 1269
rect 3708 1266 3968 1362
rect 3902 1242 3968 1266
rect 6824 1242 6834 1378
rect 3902 1237 6834 1242
rect 3902 1236 4044 1237
rect 2182 1189 2400 1213
rect 2182 1133 2302 1189
rect 2358 1133 2400 1189
rect 2182 1102 2400 1133
rect 4006 1056 6672 1064
rect 4000 1018 6672 1056
rect 4000 962 4020 1018
rect 4076 962 4100 1018
rect 4156 962 4180 1018
rect 4236 962 4260 1018
rect 4316 962 4340 1018
rect 4396 962 4420 1018
rect 4476 962 4500 1018
rect 4556 962 4580 1018
rect 4636 962 4660 1018
rect 4716 962 4740 1018
rect 4796 962 4820 1018
rect 4876 962 4900 1018
rect 4956 962 4980 1018
rect 5036 962 5060 1018
rect 5116 962 5140 1018
rect 5196 962 5220 1018
rect 5276 962 5300 1018
rect 5356 962 5380 1018
rect 5436 962 5460 1018
rect 5516 962 5540 1018
rect 5596 962 5620 1018
rect 5676 962 5700 1018
rect 5756 962 5780 1018
rect 5836 962 5860 1018
rect 5916 962 5940 1018
rect 5996 962 6020 1018
rect 6076 962 6100 1018
rect 6156 962 6180 1018
rect 6236 962 6260 1018
rect 6316 962 6340 1018
rect 6396 962 6420 1018
rect 6476 962 6500 1018
rect 6556 962 6580 1018
rect 6636 962 6672 1018
rect 4000 918 6672 962
rect 8272 1052 8580 1148
rect 4000 880 6448 918
rect 4004 860 6448 880
rect 8272 888 8590 1052
rect 8272 849 8436 888
rect 8272 793 8325 849
rect 8381 793 8436 849
rect 8272 769 8436 793
rect 8272 713 8325 769
rect 8381 713 8436 769
rect 8272 689 8436 713
rect 8272 633 8325 689
rect 8381 633 8436 689
rect 8272 556 8436 633
rect -10 208 166 243
rect -10 -16 6 208
rect 150 -16 166 208
rect 10518 213 10702 262
rect 6926 194 7020 198
rect 6918 191 7030 194
rect 6918 127 6942 191
rect 7006 127 7030 191
rect 6918 111 7030 127
rect 6918 47 6942 111
rect 7006 47 7030 111
rect 6918 44 7030 47
rect 10518 149 10572 213
rect 10636 149 10702 213
rect 10518 133 10702 149
rect 10518 69 10572 133
rect 10636 69 10702 133
rect 10518 53 10702 69
rect 6926 40 7020 44
rect -10 -51 166 -16
rect 10518 -11 10572 53
rect 10636 -11 10702 53
rect 10518 -72 10702 -11
<< via3 >>
rect 6 204 150 208
rect 6 -12 10 204
rect 10 -12 146 204
rect 146 -12 150 204
rect 6 -16 150 -12
rect 6942 127 7006 191
rect 6942 47 7006 111
rect 10572 149 10636 213
rect 10572 69 10636 133
rect 10572 -11 10636 53
<< metal4 >>
rect -15 213 10686 244
rect -15 208 10572 213
rect -15 -16 6 208
rect 150 191 10572 208
rect 150 127 6942 191
rect 7006 149 10572 191
rect 10636 149 10686 213
rect 7006 133 10686 149
rect 7006 127 10572 133
rect 150 111 10572 127
rect 150 47 6942 111
rect 7006 69 10572 111
rect 10636 69 10686 133
rect 7006 53 10686 69
rect 7006 47 10572 53
rect 150 -11 10572 47
rect 10636 -11 10686 53
rect 150 -16 10686 -11
rect -15 -54 10686 -16
use biaspmos  biaspmos_0
timestamp 1627926120
transform 1 0 4116 0 1 3370
box -52 -1706 4314 -516
use Stage2_inv  Stage2_inv_0
timestamp 1627926120
transform 1 0 2512 0 1 1150
box -102 -170 1308 1530
use Stage2_inv  Stage2_inv_1
timestamp 1627926120
transform -1 0 8210 0 1 224
box -102 -170 1308 1530
use biasnmos  biasnmos_0
timestamp 1627926120
transform 1 0 2416 0 1 90
box -70 -320 4224 814
use Stage1_inv  Stage1_inv_0
timestamp 1627926120
transform -1 0 10370 0 1 1184
box -166 -1292 1986 1598
use Stage1_inv  Stage1_inv_1
timestamp 1627926120
transform 1 0 362 0 1 1178
box -166 -1292 1986 1598
use sky130_fd_pr__res_xhigh_po_0p35_NZHUVC  sky130_fd_pr__res_xhigh_po_0p35_NZHUVC_0
timestamp 1627926120
transform 0 1 -842 -1 0 741
box -35 -508 35 508
use sky130_fd_pr__res_xhigh_po_0p35_NZHUVC  sky130_fd_pr__res_xhigh_po_0p35_NZHUVC_1
timestamp 1627926120
transform 0 1 -844 -1 0 423
box -35 -508 35 508
use sky130_fd_pr__res_xhigh_po_0p35_NZHUVC  sky130_fd_pr__res_xhigh_po_0p35_NZHUVC_2
timestamp 1627926120
transform 0 1 -840 -1 0 93
box -35 -508 35 508
<< labels >>
rlabel metal2 s 78 2790 10680 2896 4 VDD
port 1 nsew
rlabel metal2 s 110 -220 10712 -114 4 GND
port 2 nsew
rlabel metal1 s 10448 716 10622 1604 4 in2
port 3 nsew
rlabel metal1 s 126 728 222 1632 4 in1
port 4 nsew
rlabel metal1 s -748 722 100 1096 4 in
port 5 nsew
rlabel metal3 s 10526 -62 10694 254 4 out
port 6 nsew
<< end >>
