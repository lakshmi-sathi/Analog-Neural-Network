magic
tech sky130A
magscale 1 2
timestamp 1627668659
<< xpolycontact >>
rect -35 76 35 508
rect -35 -508 35 -76
<< xpolyres >>
rect -35 -76 35 76
<< viali >>
rect -19 93 19 490
rect -19 -490 19 -93
<< metal1 >>
rect -25 490 25 502
rect -25 93 -19 490
rect 19 93 25 490
rect -25 81 25 93
rect -25 -93 25 -81
rect -25 -490 -19 -93
rect 19 -490 25 -93
rect -25 -502 25 -490
<< res0p35 >>
rect -37 -78 37 78
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 0.76 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.028k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
