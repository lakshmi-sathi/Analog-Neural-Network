magic
tech sky130A
magscale 1 2
timestamp 1628045315
<< nwell >>
rect 518 1248 582 1268
rect 710 1248 774 1264
rect 902 1248 966 1266
rect 518 1222 612 1248
rect 518 1208 596 1222
rect 710 1218 804 1248
rect 902 1220 996 1248
rect 710 1208 786 1218
rect 902 1208 980 1220
rect 518 1118 582 1208
rect 710 1114 774 1208
rect 902 1116 966 1208
rect 1094 1120 1158 1270
rect 612 332 684 566
rect 604 292 684 332
rect 678 148 708 158
rect 870 148 900 158
rect 564 96 1030 148
rect 1062 142 1092 158
<< pwell >>
rect 68 768 142 1184
<< poly >>
rect 1062 105 1092 151
rect 1009 101 1092 105
rect 997 75 1092 101
<< locali >>
rect 478 1392 1194 1408
rect 478 1350 498 1392
rect 1180 1350 1194 1392
rect 478 1336 1194 1350
rect -38 -46 46 10
<< viali >>
rect 498 1350 1180 1392
<< metal1 >>
rect 482 1400 1188 1404
rect 482 1392 528 1400
rect 1146 1392 1188 1400
rect 482 1350 498 1392
rect 1180 1350 1188 1392
rect 482 1342 528 1350
rect 1146 1342 1188 1350
rect 482 1336 1188 1342
rect 128 1222 190 1276
rect 656 1202 1120 1250
rect 68 1176 142 1184
rect 68 768 76 1176
rect 128 768 142 1176
rect 518 1166 582 1174
rect 518 808 524 1166
rect 576 808 582 1166
rect 710 1166 774 1174
rect 710 828 716 1166
rect 768 828 774 1166
rect 902 1166 966 1174
rect 902 834 908 1166
rect 960 834 966 1166
rect 1094 1166 1158 1174
rect 1094 806 1100 1166
rect 1152 806 1158 1166
rect 174 164 180 556
rect 232 164 240 556
rect 614 170 620 540
rect 672 170 680 540
rect 614 164 680 170
rect 806 170 812 540
rect 864 170 872 540
rect 806 164 872 170
rect 998 170 1004 538
rect 1056 170 1064 538
rect 998 164 1064 170
rect 174 158 240 164
rect 564 120 1030 122
rect -102 32 1030 120
<< via1 >>
rect 528 1392 1146 1400
rect 528 1350 1146 1392
rect 528 1342 1146 1350
rect 76 768 128 1176
rect 524 808 576 1166
rect 716 828 768 1166
rect 908 834 960 1166
rect 1100 806 1152 1166
rect 180 164 232 556
rect 620 170 672 540
rect 812 170 864 540
rect 1004 170 1056 538
<< metal2 >>
rect -50 1426 1308 1530
rect 518 1400 1158 1426
rect 518 1342 528 1400
rect 1146 1342 1158 1400
rect 518 1262 1158 1342
rect 68 1176 142 1184
rect 68 859 76 1176
rect -25 768 76 859
rect 128 768 142 1176
rect 518 1166 582 1262
rect 518 808 524 1166
rect 576 808 582 1166
rect 710 1166 774 1262
rect 710 828 716 1166
rect 768 828 774 1166
rect 902 1166 966 1262
rect 902 834 908 1166
rect 960 834 966 1166
rect 1094 1166 1158 1262
rect 1094 806 1100 1166
rect 1152 806 1158 1166
rect -25 763 141 768
rect -25 -66 37 763
rect 174 556 240 566
rect 174 164 180 556
rect 236 172 240 556
rect 614 540 680 550
rect 232 164 240 172
rect 174 158 240 164
rect 612 174 618 540
rect 674 174 680 540
rect 612 170 620 174
rect 672 170 680 174
rect 612 160 680 170
rect 804 540 872 550
rect 804 174 810 540
rect 866 174 872 540
rect 804 170 812 174
rect 864 170 872 174
rect 804 160 872 170
rect 996 538 1064 550
rect 996 174 1002 538
rect 1058 174 1064 538
rect 996 170 1004 174
rect 1056 170 1064 174
rect 996 160 1064 170
rect -58 -170 1300 -66
<< via2 >>
rect 180 172 232 556
rect 232 172 236 556
rect 618 174 620 540
rect 620 174 672 540
rect 672 174 674 540
rect 810 174 812 540
rect 812 174 864 540
rect 864 174 866 540
rect 1002 174 1004 538
rect 1004 174 1056 538
rect 1056 174 1058 538
<< metal3 >>
rect 174 556 242 566
rect 172 304 180 556
rect 174 172 180 304
rect 236 212 250 556
rect 612 540 682 550
rect 804 540 872 550
rect 612 212 618 540
rect 236 174 618 212
rect 674 306 684 540
rect 802 306 810 540
rect 674 212 682 306
rect 804 212 810 306
rect 674 174 810 212
rect 866 212 872 540
rect 996 538 1064 550
rect 994 212 1002 538
rect 866 174 1002 212
rect 1058 350 1064 538
rect 1058 212 1068 350
rect 1058 174 1308 212
rect 236 172 1308 174
rect 174 118 1308 172
rect 174 116 1292 118
use sky130_fd_pr__nfet_01v8_LW2HKK  sky130_fd_pr__nfet_01v8_LW2HKK_0
timestamp 1627668659
transform 1 0 161 0 1 670
box -211 -730 211 730
use sky130_fd_pr__pfet_01v8_27F7GK  sky130_fd_pr__pfet_01v8_27F7GK_0
timestamp 1627668659
transform 1 0 837 0 1 661
box -455 -719 455 719
<< labels >>
rlabel metal1 -102 32 -28 120 1 in
port 3 n
rlabel metal2 -54 -164 1294 -72 1 vl
port 9 n
rlabel locali -32 -40 40 4 1 nbody
port 10 n
rlabel metal2 -44 1430 1302 1524 1 vh
port 8 n
rlabel metal3 1208 122 1304 208 1 out
port 11 n
<< end >>
