magic
tech sky130A
magscale 1 2
timestamp 1628066341
<< error_p >>
rect -269 481 -211 487
rect -77 481 -19 487
rect 115 481 173 487
rect 307 481 365 487
rect -269 447 -257 481
rect -77 447 -65 481
rect 115 447 127 481
rect 307 447 319 481
rect -269 441 -211 447
rect -77 441 -19 447
rect 115 441 173 447
rect 307 441 365 447
rect -365 -447 -307 -441
rect -173 -447 -115 -441
rect 19 -447 77 -441
rect 211 -447 269 -441
rect -365 -481 -353 -447
rect -173 -481 -161 -447
rect 19 -481 31 -447
rect 211 -481 223 -447
rect -365 -487 -307 -481
rect -173 -487 -115 -481
rect 19 -487 77 -481
rect 211 -487 269 -481
<< nwell >>
rect -551 -619 551 619
<< pmos >>
rect -351 -400 -321 400
rect -255 -400 -225 400
rect -159 -400 -129 400
rect -63 -400 -33 400
rect 33 -400 63 400
rect 129 -400 159 400
rect 225 -400 255 400
rect 321 -400 351 400
<< pdiff >>
rect -413 388 -351 400
rect -413 -388 -401 388
rect -367 -388 -351 388
rect -413 -400 -351 -388
rect -321 388 -255 400
rect -321 -388 -305 388
rect -271 -388 -255 388
rect -321 -400 -255 -388
rect -225 388 -159 400
rect -225 -388 -209 388
rect -175 -388 -159 388
rect -225 -400 -159 -388
rect -129 388 -63 400
rect -129 -388 -113 388
rect -79 -388 -63 388
rect -129 -400 -63 -388
rect -33 388 33 400
rect -33 -388 -17 388
rect 17 -388 33 388
rect -33 -400 33 -388
rect 63 388 129 400
rect 63 -388 79 388
rect 113 -388 129 388
rect 63 -400 129 -388
rect 159 388 225 400
rect 159 -388 175 388
rect 209 -388 225 388
rect 159 -400 225 -388
rect 255 388 321 400
rect 255 -388 271 388
rect 305 -388 321 388
rect 255 -400 321 -388
rect 351 388 413 400
rect 351 -388 367 388
rect 401 -388 413 388
rect 351 -400 413 -388
<< pdiffc >>
rect -401 -388 -367 388
rect -305 -388 -271 388
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect 271 -388 305 388
rect 367 -388 401 388
<< nsubdiff >>
rect -515 549 -419 583
rect 419 549 515 583
rect -515 487 -481 549
rect 481 487 515 549
rect -515 -549 -481 -487
rect 481 -549 515 -487
rect -515 -583 -419 -549
rect 419 -583 515 -549
<< nsubdiffcont >>
rect -419 549 419 583
rect -515 -487 -481 487
rect 481 -487 515 487
rect -419 -583 419 -549
<< poly >>
rect -273 481 -207 497
rect -273 447 -257 481
rect -223 447 -207 481
rect -273 431 -207 447
rect -81 481 -15 497
rect -81 447 -65 481
rect -31 447 -15 481
rect -81 431 -15 447
rect 111 481 177 497
rect 111 447 127 481
rect 161 447 177 481
rect 111 431 177 447
rect 303 481 369 497
rect 303 447 319 481
rect 353 447 369 481
rect 303 431 369 447
rect -351 400 -321 426
rect -255 400 -225 431
rect -159 400 -129 426
rect -63 400 -33 431
rect 33 400 63 426
rect 129 400 159 431
rect 225 400 255 426
rect 321 400 351 431
rect -351 -431 -321 -400
rect -255 -426 -225 -400
rect -159 -431 -129 -400
rect -63 -426 -33 -400
rect 33 -431 63 -400
rect 129 -426 159 -400
rect 225 -431 255 -400
rect 321 -426 351 -400
rect -369 -447 -303 -431
rect -369 -481 -353 -447
rect -319 -481 -303 -447
rect -369 -497 -303 -481
rect -177 -447 -111 -431
rect -177 -481 -161 -447
rect -127 -481 -111 -447
rect -177 -497 -111 -481
rect 15 -447 81 -431
rect 15 -481 31 -447
rect 65 -481 81 -447
rect 15 -497 81 -481
rect 207 -447 273 -431
rect 207 -481 223 -447
rect 257 -481 273 -447
rect 207 -497 273 -481
<< polycont >>
rect -257 447 -223 481
rect -65 447 -31 481
rect 127 447 161 481
rect 319 447 353 481
rect -353 -481 -319 -447
rect -161 -481 -127 -447
rect 31 -481 65 -447
rect 223 -481 257 -447
<< locali >>
rect -515 549 -419 583
rect 419 549 515 583
rect -515 487 -481 549
rect 481 487 515 549
rect -273 447 -257 481
rect -223 447 -207 481
rect -81 447 -65 481
rect -31 447 -15 481
rect 111 447 127 481
rect 161 447 177 481
rect 303 447 319 481
rect 353 447 369 481
rect -401 388 -367 404
rect -401 -404 -367 -388
rect -305 388 -271 404
rect -305 -404 -271 -388
rect -209 388 -175 404
rect -209 -404 -175 -388
rect -113 388 -79 404
rect -113 -404 -79 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 79 388 113 404
rect 79 -404 113 -388
rect 175 388 209 404
rect 175 -404 209 -388
rect 271 388 305 404
rect 271 -404 305 -388
rect 367 388 401 404
rect 367 -404 401 -388
rect -369 -481 -353 -447
rect -319 -481 -303 -447
rect -177 -481 -161 -447
rect -127 -481 -111 -447
rect 15 -481 31 -447
rect 65 -481 81 -447
rect 207 -481 223 -447
rect 257 -481 273 -447
rect -515 -549 -481 -487
rect 481 -549 515 -487
rect -515 -583 -419 -549
rect 419 -583 515 -549
<< viali >>
rect -257 447 -223 481
rect -65 447 -31 481
rect 127 447 161 481
rect 319 447 353 481
rect -401 -388 -367 388
rect -305 -388 -271 388
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect 271 -388 305 388
rect 367 -388 401 388
rect -353 -481 -319 -447
rect -161 -481 -127 -447
rect 31 -481 65 -447
rect 223 -481 257 -447
<< metal1 >>
rect -269 481 -211 487
rect -269 447 -257 481
rect -223 447 -211 481
rect -269 441 -211 447
rect -77 481 -19 487
rect -77 447 -65 481
rect -31 447 -19 481
rect -77 441 -19 447
rect 115 481 173 487
rect 115 447 127 481
rect 161 447 173 481
rect 115 441 173 447
rect 307 481 365 487
rect 307 447 319 481
rect 353 447 365 481
rect 307 441 365 447
rect -407 388 -361 400
rect -407 -388 -401 388
rect -367 -388 -361 388
rect -407 -400 -361 -388
rect -311 388 -265 400
rect -311 -388 -305 388
rect -271 -388 -265 388
rect -311 -400 -265 -388
rect -215 388 -169 400
rect -215 -388 -209 388
rect -175 -388 -169 388
rect -215 -400 -169 -388
rect -119 388 -73 400
rect -119 -388 -113 388
rect -79 -388 -73 388
rect -119 -400 -73 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 73 388 119 400
rect 73 -388 79 388
rect 113 -388 119 388
rect 73 -400 119 -388
rect 169 388 215 400
rect 169 -388 175 388
rect 209 -388 215 388
rect 169 -400 215 -388
rect 265 388 311 400
rect 265 -388 271 388
rect 305 -388 311 388
rect 265 -400 311 -388
rect 361 388 407 400
rect 361 -388 367 388
rect 401 -388 407 388
rect 361 -400 407 -388
rect -365 -447 -307 -441
rect -365 -481 -353 -447
rect -319 -481 -307 -447
rect -365 -487 -307 -481
rect -173 -447 -115 -441
rect -173 -481 -161 -447
rect -127 -481 -115 -447
rect -173 -487 -115 -481
rect 19 -447 77 -441
rect 19 -481 31 -447
rect 65 -481 77 -447
rect 19 -487 77 -481
rect 211 -447 269 -441
rect 211 -481 223 -447
rect 257 -481 269 -447
rect 211 -487 269 -481
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -498 -566 498 566
string parameters w 4 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
