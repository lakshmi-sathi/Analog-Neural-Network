magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_s >>
rect 15088 4915 15446 4984
rect 15256 4816 15278 4915
rect 15352 4816 15446 4915
rect 49774 4913 50132 4982
rect 84028 4917 84386 4986
rect 15256 4815 15446 4816
rect 15220 4709 15446 4815
rect 49942 4814 49964 4913
rect 50038 4814 50132 4913
rect 84196 4818 84218 4917
rect 84292 4818 84386 4917
rect 84196 4817 84386 4818
rect 49942 4813 50132 4814
rect 15220 4671 15314 4709
rect 15352 4671 15446 4709
rect 15220 4647 15446 4671
rect 49906 4707 50132 4813
rect 49906 4669 50000 4707
rect 50038 4669 50132 4707
rect 49906 4645 50132 4669
rect 84160 4711 84386 4817
rect 84160 4673 84254 4711
rect 84292 4673 84386 4711
rect 84160 4649 84386 4673
rect 15096 3661 15454 3730
rect 15264 3562 15286 3661
rect 15360 3562 15454 3661
rect 49782 3659 50140 3728
rect 84036 3663 84394 3732
rect 15264 3561 15454 3562
rect 15228 3455 15454 3561
rect 49950 3560 49972 3659
rect 50046 3560 50140 3659
rect 84204 3564 84226 3663
rect 84300 3564 84394 3663
rect 84204 3563 84394 3564
rect 49950 3559 50140 3560
rect 15228 3417 15322 3455
rect 15360 3417 15454 3455
rect 15228 3393 15454 3417
rect 49914 3453 50140 3559
rect 49914 3415 50008 3453
rect 50046 3415 50140 3453
rect 49914 3391 50140 3415
rect 84168 3457 84394 3563
rect 84168 3419 84262 3457
rect 84300 3419 84394 3457
rect 84168 3395 84394 3419
rect 15076 2393 15434 2462
rect 15244 2294 15266 2393
rect 15340 2294 15434 2393
rect 49762 2391 50120 2460
rect 84016 2395 84374 2464
rect 15244 2293 15434 2294
rect 15208 2187 15434 2293
rect 49930 2292 49952 2391
rect 50026 2292 50120 2391
rect 84184 2296 84206 2395
rect 84280 2296 84374 2395
rect 84184 2295 84374 2296
rect 49930 2291 50120 2292
rect 15208 2149 15302 2187
rect 15340 2149 15434 2187
rect 15208 2125 15434 2149
rect 49894 2185 50120 2291
rect 49894 2147 49988 2185
rect 50026 2147 50120 2185
rect 49894 2123 50120 2147
rect 84148 2189 84374 2295
rect 84148 2151 84242 2189
rect 84280 2151 84374 2189
rect 84148 2127 84374 2151
rect 15078 -2106 15436 -2000
rect 15246 -2168 15268 -2106
rect 15342 -2168 15436 -2106
rect 49764 -2108 50122 -2002
rect 84018 -2104 84376 -1998
rect 15210 -2192 15436 -2168
rect 49932 -2170 49954 -2108
rect 50028 -2170 50122 -2108
rect 84186 -2166 84208 -2104
rect 84282 -2166 84376 -2104
rect 15210 -2230 15304 -2192
rect 15342 -2230 15436 -2192
rect 15210 -2336 15436 -2230
rect 15246 -2337 15436 -2336
rect 49896 -2194 50122 -2170
rect 49896 -2232 49990 -2194
rect 50028 -2232 50122 -2194
rect 49896 -2338 50122 -2232
rect 84150 -2190 84376 -2166
rect 84150 -2228 84244 -2190
rect 84282 -2228 84376 -2190
rect 84150 -2334 84376 -2228
rect 84186 -2335 84376 -2334
rect 49932 -2339 50122 -2338
rect 15098 -3374 15456 -3268
rect 15266 -3436 15288 -3374
rect 15362 -3436 15456 -3374
rect 49784 -3376 50142 -3270
rect 84038 -3372 84396 -3266
rect 15230 -3460 15456 -3436
rect 49952 -3438 49974 -3376
rect 50048 -3438 50142 -3376
rect 84206 -3434 84228 -3372
rect 84302 -3434 84396 -3372
rect 15230 -3498 15324 -3460
rect 15362 -3498 15456 -3460
rect 15230 -3604 15456 -3498
rect 15266 -3605 15456 -3604
rect 49916 -3462 50142 -3438
rect 49916 -3500 50010 -3462
rect 50048 -3500 50142 -3462
rect 49916 -3606 50142 -3500
rect 84170 -3458 84396 -3434
rect 84170 -3496 84264 -3458
rect 84302 -3496 84396 -3458
rect 84170 -3602 84396 -3496
rect 84206 -3603 84396 -3602
rect 49952 -3607 50142 -3606
rect 15090 -4628 15448 -4522
rect 15258 -4690 15280 -4628
rect 15354 -4690 15448 -4628
rect 49776 -4630 50134 -4524
rect 84030 -4626 84388 -4520
rect 15222 -4714 15448 -4690
rect 49944 -4692 49966 -4630
rect 50040 -4692 50134 -4630
rect 84198 -4688 84220 -4626
rect 84294 -4688 84388 -4626
rect 15222 -4752 15316 -4714
rect 15354 -4752 15448 -4714
rect 15222 -4858 15448 -4752
rect 15258 -4859 15448 -4858
rect 49908 -4716 50134 -4692
rect 49908 -4754 50002 -4716
rect 50040 -4754 50134 -4716
rect 49908 -4860 50134 -4754
rect 84162 -4712 84388 -4688
rect 84162 -4750 84256 -4712
rect 84294 -4750 84388 -4712
rect 84162 -4856 84388 -4750
rect 84198 -4857 84388 -4856
rect 49944 -4861 50134 -4860
rect 15000 -14011 15358 -13942
rect 15168 -14110 15190 -14011
rect 15264 -14110 15358 -14011
rect 49686 -14013 50044 -13944
rect 15168 -14111 15358 -14110
rect 15132 -14217 15358 -14111
rect 49854 -14112 49876 -14013
rect 49950 -14112 50044 -14013
rect 49854 -14113 50044 -14112
rect 15132 -14255 15226 -14217
rect 15264 -14255 15358 -14217
rect 15132 -14279 15358 -14255
rect 49818 -14219 50044 -14113
rect 49818 -14257 49912 -14219
rect 49950 -14257 50044 -14219
rect 49818 -14281 50044 -14257
rect 15008 -15265 15366 -15196
rect 15176 -15364 15198 -15265
rect 15272 -15364 15366 -15265
rect 49694 -15267 50052 -15198
rect 15176 -15365 15366 -15364
rect 15140 -15471 15366 -15365
rect 49862 -15366 49884 -15267
rect 49958 -15366 50052 -15267
rect 49862 -15367 50052 -15366
rect 15140 -15509 15234 -15471
rect 15272 -15509 15366 -15471
rect 15140 -15533 15366 -15509
rect 49826 -15473 50052 -15367
rect 49826 -15511 49920 -15473
rect 49958 -15511 50052 -15473
rect 49826 -15535 50052 -15511
rect 14988 -16533 15346 -16464
rect 15156 -16632 15178 -16533
rect 15252 -16632 15346 -16533
rect 49674 -16535 50032 -16466
rect 15156 -16633 15346 -16632
rect 15120 -16739 15346 -16633
rect 49842 -16634 49864 -16535
rect 49938 -16634 50032 -16535
rect 49842 -16635 50032 -16634
rect 15120 -16777 15214 -16739
rect 15252 -16777 15346 -16739
rect 15120 -16801 15346 -16777
rect 49806 -16741 50032 -16635
rect 49806 -16779 49900 -16741
rect 49938 -16779 50032 -16741
rect 49806 -16803 50032 -16779
<< locali >>
rect 14006 6337 14226 6358
rect 14006 6159 14027 6337
rect 14205 6159 14226 6337
rect 14006 3816 14226 6159
rect 49509 5293 50017 5304
rect 14821 5240 15334 5262
rect 14821 5134 15206 5240
rect 15312 5134 15334 5240
rect 14821 5113 15334 5134
rect 49509 5187 49900 5293
rect 50006 5187 50017 5293
rect 49509 5177 50017 5187
rect 83736 5274 84284 5304
rect 14821 4973 14968 5113
rect 49509 4971 49654 5177
rect 83736 5168 84148 5274
rect 84254 5168 84284 5274
rect 83736 5139 84284 5168
rect 83736 4975 83908 5139
rect 14006 3719 14733 3816
rect 14014 2548 14229 3719
rect 49490 2655 49987 2668
rect 49490 2549 49868 2655
rect 49974 2549 49987 2655
rect 14014 2451 14856 2548
rect 49490 2537 49987 2549
rect 49490 2449 49639 2537
rect 82825 2453 83682 2550
rect 82825 279 83070 2453
rect 82825 101 82858 279
rect 83036 101 83070 279
rect 82825 68 83070 101
rect 82912 32 83070 68
rect 13888 -12578 14063 -12543
rect 13888 -12684 13922 -12578
rect 14028 -12684 14063 -12578
rect 13888 -15110 14063 -12684
rect 49257 -12599 49475 -12579
rect 49257 -12777 49277 -12599
rect 49455 -12777 49475 -12599
rect 49257 -13335 49475 -12777
rect 14716 -13597 15246 -13578
rect 14716 -13703 15114 -13597
rect 15220 -13671 15246 -13597
rect 48563 -13599 49475 -13335
rect 15220 -13703 15239 -13671
rect 14716 -13721 15239 -13703
rect 14716 -13952 14870 -13721
rect 13888 -15207 14714 -15110
rect 13894 -16378 14070 -15207
rect 13894 -16475 14697 -16378
rect 48563 -16380 48781 -13599
rect 49257 -13954 49475 -13599
rect 48563 -16457 49499 -16380
rect 48606 -16477 49499 -16457
<< viali >>
rect 14027 6159 14205 6337
rect 15206 5134 15312 5240
rect 49900 5187 50006 5293
rect 84148 5168 84254 5274
rect 49868 2549 49974 2655
rect 82858 101 83036 279
rect 13922 -12684 14028 -12578
rect 49277 -12777 49455 -12599
rect 15114 -13703 15220 -13597
<< metal1 >>
rect 34608 8319 35192 8322
rect 34 8184 464 8190
rect 34 7684 63 8184
rect 435 7684 464 8184
rect 34 7678 464 7684
rect 34608 7627 34618 8319
rect 35182 7627 35192 8319
rect 68926 8256 69410 8292
rect 68926 7756 68993 8256
rect 69365 7756 69410 8256
rect 68926 7664 69410 7756
rect 34608 7624 35192 7627
rect 13994 6338 14238 6364
rect 13994 6158 14026 6338
rect 14206 6158 14238 6338
rect 13994 6132 14238 6158
rect 49878 5298 50029 5310
rect 15173 5245 15346 5268
rect 15173 5129 15201 5245
rect 15317 5129 15346 5245
rect 49878 5182 49895 5298
rect 50011 5182 50029 5298
rect 49878 5171 50029 5182
rect 84107 5279 84296 5310
rect 84107 5163 84143 5279
rect 84259 5163 84296 5279
rect 84107 5133 84296 5163
rect 15173 5107 15346 5129
rect 34714 4732 35132 4734
rect 18 4701 454 4726
rect 18 4265 50 4701
rect 422 4265 454 4701
rect 15530 4476 16376 4696
rect 18092 4468 18964 4704
rect 18 4240 454 4265
rect 34714 4232 34737 4732
rect 35109 4232 35132 4732
rect 68966 4712 69424 4738
rect 50208 4477 51353 4699
rect 52204 4474 53756 4698
rect 68966 4276 68977 4712
rect 69413 4276 69424 4712
rect 84450 4481 85479 4703
rect 86807 4480 87980 4702
rect 68966 4250 69424 4276
rect 34714 4230 35132 4232
rect 15546 3244 16942 3456
rect 17249 3276 19040 3498
rect 49844 2660 49999 2674
rect 49844 2544 49863 2660
rect 49979 2544 49999 2660
rect 49844 2531 49999 2544
rect 15509 1986 16941 2188
rect 17583 2000 19038 2218
rect 50234 1984 51497 2186
rect 52279 1998 53724 2216
rect 84488 1988 85859 2190
rect 86479 2002 87978 2220
rect 32527 1938 35228 1958
rect 28 1909 480 1930
rect 28 1473 68 1909
rect 440 1473 480 1909
rect 28 1452 480 1473
rect 32527 1438 32554 1938
rect 32990 1438 35228 1938
rect 32527 1416 35228 1438
rect 66955 1915 69781 1962
rect 66955 1479 67053 1915
rect 67489 1479 69781 1915
rect 66955 1420 69781 1479
rect 82813 312 83082 319
rect 82813 68 82825 312
rect 83069 68 83082 312
rect 82813 62 83082 68
rect 46 -1485 514 -1484
rect 46 -1985 62 -1485
rect 498 -1985 514 -1485
rect 46 -1986 514 -1985
rect 32513 -1488 35230 -1463
rect 32513 -1988 32572 -1488
rect 33008 -1988 35230 -1488
rect 68976 -1516 69414 -1496
rect 68976 -1952 69009 -1516
rect 69381 -1952 69414 -1516
rect 68976 -1972 69414 -1952
rect 32513 -2005 35230 -1988
rect 18920 -2178 20268 -2146
rect 18920 -3254 19546 -2178
rect 20174 -2346 20268 -2178
rect 84490 -2229 85755 -2027
rect 53606 -2274 54968 -2232
rect 86395 -2259 87980 -2041
rect 20174 -2706 20290 -2346
rect 20174 -3254 20281 -2706
rect 18920 -3270 20281 -3254
rect 53606 -3222 54151 -2274
rect 54907 -2832 54968 -2274
rect 54907 -2910 54952 -2832
rect 54907 -3222 54962 -2910
rect 53606 -3270 54962 -3222
rect 19508 -3280 20212 -3270
rect 20 -4342 450 -4324
rect 20 -4778 49 -4342
rect 421 -4778 450 -4342
rect 20 -4796 450 -4778
rect 34726 -4331 35046 -4302
rect 34726 -4767 34764 -4331
rect 35008 -4767 35046 -4331
rect 34726 -4796 35046 -4767
rect 68976 -4322 69434 -4296
rect 68976 -4758 68987 -4322
rect 69423 -4758 69434 -4322
rect 68976 -4784 69434 -4758
rect 72 -7731 442 -7728
rect 72 -8231 103 -7731
rect 411 -8231 442 -7731
rect 66961 -7733 69573 -7709
rect 72 -8234 442 -8231
rect 34730 -7781 35136 -7758
rect 34730 -8217 34747 -7781
rect 35119 -8217 35136 -7781
rect 34730 -8240 35136 -8217
rect 66961 -8233 67005 -7733
rect 67505 -8233 69573 -7733
rect 66961 -8251 69573 -8233
rect -32 -10765 354 -10754
rect -32 -11201 7 -10765
rect 315 -11201 354 -10765
rect -32 -11212 354 -11201
rect 34642 -10794 35056 -10764
rect 34642 -11230 34663 -10794
rect 35035 -11230 35056 -10794
rect 34642 -11260 35056 -11230
rect 13876 -12573 14075 -12537
rect 13876 -12689 13917 -12573
rect 14033 -12689 14075 -12573
rect 13876 -12724 14075 -12689
rect 49245 -12598 49487 -12573
rect 49245 -12778 49276 -12598
rect 49456 -12778 49487 -12598
rect 49245 -12803 49487 -12778
rect 15084 -13592 15251 -13572
rect 15084 -13708 15109 -13592
rect 15225 -13708 15251 -13592
rect 15084 -13727 15251 -13708
rect -58 -14181 304 -14180
rect -58 -14681 -31 -14181
rect 277 -14681 304 -14181
rect 34632 -14214 35036 -14192
rect 15434 -14447 16271 -14225
rect 18100 -14450 18982 -14226
rect 34632 -14650 34648 -14214
rect 35020 -14650 35036 -14214
rect 50120 -14449 51119 -14227
rect 52490 -14452 53668 -14228
rect 34632 -14672 35036 -14650
rect -58 -14682 304 -14681
rect 15432 -15682 16914 -15470
rect 17237 -15650 18952 -15428
rect 15437 -16940 16881 -16738
rect 17439 -16926 18950 -16708
rect 50146 -16942 50962 -16740
rect 52121 -16928 53636 -16710
rect -80 -16985 320 -16974
rect -80 -17485 -66 -16985
rect 306 -17485 320 -16985
rect -80 -17496 320 -17485
rect 34598 -17000 35056 -16998
rect 34598 -17500 34609 -17000
rect 35045 -17500 35056 -17000
rect 34598 -17502 35056 -17500
<< via1 >>
rect 63 7684 435 8184
rect 34618 7627 35182 8319
rect 68993 7756 69365 8256
rect 14026 6337 14206 6338
rect 14026 6159 14027 6337
rect 14027 6159 14205 6337
rect 14205 6159 14206 6337
rect 14026 6158 14206 6159
rect 15201 5240 15317 5245
rect 15201 5134 15206 5240
rect 15206 5134 15312 5240
rect 15312 5134 15317 5240
rect 15201 5129 15317 5134
rect 49895 5293 50011 5298
rect 49895 5187 49900 5293
rect 49900 5187 50006 5293
rect 50006 5187 50011 5293
rect 49895 5182 50011 5187
rect 84143 5274 84259 5279
rect 84143 5168 84148 5274
rect 84148 5168 84254 5274
rect 84254 5168 84259 5274
rect 84143 5163 84259 5168
rect 50 4265 422 4701
rect 34737 4232 35109 4732
rect 68977 4276 69413 4712
rect 49863 2655 49979 2660
rect 49863 2549 49868 2655
rect 49868 2549 49974 2655
rect 49974 2549 49979 2655
rect 49863 2544 49979 2549
rect 68 1473 440 1909
rect 32554 1438 32990 1938
rect 67053 1479 67489 1915
rect 82825 279 83069 312
rect 82825 101 82858 279
rect 82858 101 83036 279
rect 83036 101 83069 279
rect 82825 68 83069 101
rect 62 -1985 498 -1485
rect 32572 -1988 33008 -1488
rect 69009 -1952 69381 -1516
rect 19546 -3254 20174 -2178
rect 54151 -3222 54907 -2274
rect 49 -4778 421 -4342
rect 34764 -4767 35008 -4331
rect 68987 -4758 69423 -4322
rect 103 -8231 411 -7731
rect 34747 -8217 35119 -7781
rect 67005 -8233 67505 -7733
rect 7 -11201 315 -10765
rect 34663 -11230 35035 -10794
rect 13917 -12578 14033 -12573
rect 13917 -12684 13922 -12578
rect 13922 -12684 14028 -12578
rect 14028 -12684 14033 -12578
rect 13917 -12689 14033 -12684
rect 49276 -12599 49456 -12598
rect 49276 -12777 49277 -12599
rect 49277 -12777 49455 -12599
rect 49455 -12777 49456 -12599
rect 49276 -12778 49456 -12777
rect 15109 -13597 15225 -13592
rect 15109 -13703 15114 -13597
rect 15114 -13703 15220 -13597
rect 15220 -13703 15225 -13597
rect 15109 -13708 15225 -13703
rect -31 -14681 277 -14181
rect 34648 -14650 35020 -14214
rect -66 -17485 306 -16985
rect 34609 -17500 35045 -17000
<< metal2 >>
rect 1460 9280 99566 9417
rect 34618 8321 35182 8332
rect 34618 8319 34632 8321
rect 35168 8319 35182 8321
rect 44 8184 454 8200
rect 44 8162 63 8184
rect 435 8162 454 8184
rect 44 7706 61 8162
rect 437 7706 454 8162
rect 44 7684 63 7706
rect 435 7684 454 7706
rect 44 7668 454 7684
rect 68962 8274 69396 8292
rect 68962 7738 68991 8274
rect 69367 7738 69396 8274
rect 68962 7720 69396 7738
rect 34618 7625 34632 7627
rect 35168 7625 35182 7627
rect 34618 7614 35182 7625
rect 14006 6338 14226 6368
rect 14006 6158 14026 6338
rect 14206 6158 14226 6338
rect 14006 6128 14226 6158
rect 64882 5856 65228 5876
rect 30222 5805 30564 5854
rect 15256 5327 15338 5677
rect 30222 5589 30245 5805
rect 30541 5589 30564 5805
rect 30222 5540 30564 5589
rect 64882 5560 64907 5856
rect 65203 5560 65228 5856
rect 64882 5540 65228 5560
rect 49890 5298 50017 5314
rect 15185 5245 15334 5272
rect 15185 5129 15201 5245
rect 15317 5129 15334 5245
rect 49890 5182 49895 5298
rect 50011 5182 50017 5298
rect 49890 5167 50017 5182
rect 84119 5279 84284 5314
rect 84119 5163 84143 5279
rect 84259 5163 84284 5279
rect 84119 5129 84284 5163
rect 15185 5103 15334 5129
rect 28 4711 444 4736
rect 28 4255 48 4711
rect 424 4255 444 4711
rect 28 4230 444 4255
rect 34724 4732 35122 4744
rect 34724 4710 34737 4732
rect 35109 4710 35122 4732
rect 34724 4254 34735 4710
rect 35111 4254 35122 4710
rect 34724 4232 34737 4254
rect 35109 4232 35122 4254
rect 68976 4722 69414 4748
rect 68976 4712 69007 4722
rect 69383 4712 69414 4722
rect 68976 4276 68977 4712
rect 69413 4276 69414 4712
rect 68976 4266 69007 4276
rect 69383 4266 69414 4276
rect 68976 4240 69414 4266
rect 34724 4220 35122 4232
rect 49856 2660 49987 2678
rect 49856 2544 49863 2660
rect 49979 2544 49987 2660
rect 49856 2527 49987 2544
rect -8550 1427 -7096 2048
rect -5372 1938 -4186 1953
rect 38 1938 470 1940
rect -5382 1909 470 1938
rect -5382 1480 68 1909
rect -8550 -69 -8337 1427
rect -7321 -69 -7096 1427
rect -8550 -546 -7096 -69
rect -5372 -1484 -4186 1480
rect 38 1473 68 1480
rect 440 1473 470 1909
rect 38 1442 470 1473
rect 32552 1938 32992 1962
rect 32552 1438 32554 1938
rect 32990 1438 32992 1938
rect 67046 1915 67496 1928
rect 67046 1479 67053 1915
rect 67489 1479 67496 1915
rect 67046 1466 67496 1479
rect 32552 1414 32992 1438
rect 82825 312 83070 323
rect 28944 238 28966 240
rect 28944 120 28974 238
rect 2022 35 19190 110
rect 2022 -150 13690 35
rect 14226 -150 19190 35
rect 21204 94 28986 120
rect 63638 100 63664 294
rect 21204 -38 54118 94
rect 21204 -140 48495 -38
rect 28658 -156 48495 -140
rect 13690 -212 14226 -181
rect 28944 -268 28974 -156
rect 28946 -274 28974 -268
rect 48456 -254 48495 -156
rect 48951 -156 54118 -38
rect 55562 68 82825 100
rect 83069 100 83070 312
rect 97884 124 97912 242
rect 83069 68 88342 100
rect 48951 -254 48992 -156
rect 55562 -162 88342 68
rect 48456 -288 48992 -254
rect 63638 -276 63664 -162
rect 89808 -170 97912 124
rect 97884 -282 97912 -170
rect 56 -1484 504 -1474
rect -5372 -1485 504 -1484
rect -5372 -1958 62 -1485
rect -8612 -5489 -7158 -4846
rect -8612 -6985 -8394 -5489
rect -7298 -6985 -7158 -5489
rect -8612 -7440 -7158 -6985
rect -8550 -11908 -7096 -11172
rect -5372 -11908 -4186 -1958
rect 56 -1985 62 -1958
rect 498 -1985 504 -1485
rect 56 -1996 504 -1985
rect 32570 -1488 33010 -1464
rect 32570 -1988 32572 -1488
rect 33008 -1988 33010 -1488
rect 68986 -1506 69404 -1486
rect 68986 -1962 69007 -1506
rect 69383 -1962 69404 -1506
rect 68986 -1982 69404 -1962
rect 32570 -2012 33010 -1988
rect 19518 -2178 20202 -2142
rect 19518 -3254 19546 -2178
rect 20174 -3254 20202 -2178
rect 54128 -2274 54930 -2254
rect 54128 -3222 54151 -2274
rect 54907 -3222 54930 -2274
rect 54128 -3242 54930 -3222
rect 19518 -3290 20202 -3254
rect 30 -4332 440 -4314
rect 30 -4788 47 -4332
rect 423 -4788 440 -4332
rect 30 -4806 440 -4788
rect 34736 -4321 35036 -4292
rect 34736 -4777 34738 -4321
rect 35034 -4777 35036 -4321
rect 34736 -4806 35036 -4777
rect 68986 -4312 69424 -4286
rect 68986 -4322 69017 -4312
rect 69393 -4322 69424 -4312
rect 68986 -4758 68987 -4322
rect 69423 -4758 69424 -4322
rect 68986 -4768 69017 -4758
rect 69393 -4768 69424 -4758
rect 68986 -4794 69424 -4768
rect 30208 -5590 30568 -5570
rect 30208 -5886 30240 -5590
rect 30536 -5886 30568 -5590
rect 30208 -5906 30568 -5886
rect 64870 -5616 65252 -5574
rect 64870 -5992 64873 -5616
rect 65249 -5992 65252 -5616
rect 64870 -6034 65252 -5992
rect 99112 -6733 99518 6411
rect 82 -7731 432 -7718
rect 82 -8231 103 -7731
rect 411 -8231 432 -7731
rect 66992 -7733 67518 -7714
rect 82 -8244 432 -8231
rect 34740 -7771 35126 -7748
rect 34740 -8227 34745 -7771
rect 35121 -8227 35126 -7771
rect 34740 -8250 35126 -8227
rect 66992 -8233 67005 -7733
rect 67505 -8233 67518 -7733
rect 66992 -8252 67518 -8233
rect 644 -9344 1786 -9338
rect 644 -9604 1778 -9344
rect 4370 -9378 30488 -9338
rect 4370 -9600 36660 -9378
rect 4362 -9604 36660 -9600
rect 28836 -9628 36660 -9604
rect 38876 -9628 99490 -9378
rect -22 -10755 344 -10744
rect -22 -10765 13 -10755
rect 309 -10765 344 -10755
rect -22 -11201 7 -10765
rect 315 -11201 344 -10765
rect -22 -11211 13 -11201
rect 309 -11211 344 -11201
rect -22 -11222 344 -11211
rect 34652 -10784 35046 -10754
rect 34652 -11240 34661 -10784
rect 35037 -11240 35046 -10784
rect 34652 -11270 35046 -11240
rect -8550 -13094 -4186 -11908
rect 13888 -12573 14063 -12533
rect 13888 -12689 13917 -12573
rect 14033 -12689 14063 -12573
rect 13888 -12728 14063 -12689
rect 49257 -12598 49475 -12569
rect 49257 -12778 49276 -12598
rect 49456 -12778 49475 -12598
rect 49257 -12807 49475 -12778
rect -8550 -13126 -6654 -13094
rect -8550 -13766 -7096 -13126
rect -5372 -16978 -4186 -13094
rect 15096 -13592 15239 -13568
rect 15096 -13708 15109 -13592
rect 15225 -13708 15239 -13592
rect 15096 -13731 15239 -13708
rect -48 -14181 294 -14170
rect -48 -14681 -31 -14181
rect 277 -14681 294 -14181
rect -48 -14692 294 -14681
rect 34642 -14204 35026 -14182
rect 34642 -14660 34646 -14204
rect 35022 -14660 35026 -14204
rect 34642 -14682 35026 -14660
rect -70 -16978 310 -16964
rect -5372 -16985 310 -16978
rect -5372 -17476 -66 -16985
rect -5372 -17661 -4186 -17476
rect -70 -17485 -66 -17476
rect 306 -17485 310 -16985
rect -70 -17506 310 -17485
rect 34608 -17000 35046 -16988
rect 34608 -17500 34609 -17000
rect 35045 -17500 35046 -17000
rect 34608 -17512 35046 -17500
rect 48434 -18633 49004 -18582
rect 13674 -18735 14250 -18686
rect 13674 -18808 13694 -18735
rect 2038 -18871 13694 -18808
rect 14230 -18808 14250 -18735
rect 48434 -18808 48531 -18633
rect 14230 -18849 48531 -18808
rect 48907 -18808 49004 -18633
rect 48907 -18849 63550 -18808
rect 14230 -18871 63550 -18849
rect 2038 -18920 63550 -18871
<< via2 >>
rect 34632 8319 35168 8321
rect 61 7706 63 8162
rect 63 7706 435 8162
rect 435 7706 437 8162
rect 34632 7627 35168 8319
rect 68991 8256 69367 8274
rect 68991 7756 68993 8256
rect 68993 7756 69365 8256
rect 69365 7756 69367 8256
rect 68991 7738 69367 7756
rect 34632 7625 35168 7627
rect 30245 5589 30541 5805
rect 64907 5560 65203 5856
rect 48 4701 424 4711
rect 48 4265 50 4701
rect 50 4265 422 4701
rect 422 4265 424 4701
rect 48 4255 424 4265
rect 34735 4254 34737 4710
rect 34737 4254 35109 4710
rect 35109 4254 35111 4710
rect 69007 4712 69383 4722
rect 69007 4276 69383 4712
rect 69007 4266 69383 4276
rect -8337 -69 -7321 1427
rect 32584 1460 32960 1916
rect 67083 1509 67459 1885
rect 13690 -181 14226 35
rect 48495 -254 48951 -38
rect -8394 -6985 -7298 -5489
rect 32602 -1966 32978 -1510
rect 69007 -1516 69383 -1506
rect 69007 -1952 69009 -1516
rect 69009 -1952 69381 -1516
rect 69381 -1952 69383 -1516
rect 69007 -1962 69383 -1952
rect 47 -4342 423 -4332
rect 47 -4778 49 -4342
rect 49 -4778 421 -4342
rect 421 -4778 423 -4342
rect 47 -4788 423 -4778
rect 34738 -4331 35034 -4321
rect 34738 -4767 34764 -4331
rect 34764 -4767 35008 -4331
rect 35008 -4767 35034 -4331
rect 34738 -4777 35034 -4767
rect 69017 -4322 69393 -4312
rect 69017 -4758 69393 -4322
rect 69017 -4768 69393 -4758
rect 30240 -5886 30536 -5590
rect 64873 -5992 65249 -5616
rect 109 -8209 405 -7753
rect 34745 -7781 35121 -7771
rect 34745 -8217 34747 -7781
rect 34747 -8217 35119 -7781
rect 35119 -8217 35121 -7781
rect 34745 -8227 35121 -8217
rect 67027 -8211 67483 -7755
rect 13 -10765 309 -10755
rect 13 -11201 309 -10765
rect 13 -11211 309 -11201
rect 34661 -10794 35037 -10784
rect 34661 -11230 34663 -10794
rect 34663 -11230 35035 -10794
rect 35035 -11230 35037 -10794
rect 34661 -11240 35037 -11230
rect -25 -14659 271 -14203
rect 34646 -14214 35022 -14204
rect 34646 -14650 34648 -14214
rect 34648 -14650 35020 -14214
rect 35020 -14650 35022 -14214
rect 34646 -14660 35022 -14650
rect 34639 -17478 35015 -17022
rect 13694 -18871 14230 -18735
rect 48531 -18849 48907 -18633
<< metal3 >>
rect 34608 8321 35192 8327
rect 34608 8285 34632 8321
rect 35168 8285 35192 8321
rect 34 8166 464 8195
rect 34 7702 57 8166
rect 441 7702 464 8166
rect 34 7673 464 7702
rect 34608 7661 34628 8285
rect 35172 7661 35192 8285
rect 68952 8278 69406 8287
rect 68952 7734 68987 8278
rect 69371 7734 69406 8278
rect 68952 7725 69406 7734
rect 34608 7625 34632 7661
rect 35168 7625 35192 7661
rect 34608 7619 35192 7625
rect 64872 5869 65238 5871
rect 30208 5849 30564 5862
rect 64870 5856 65252 5869
rect 30208 5805 30574 5849
rect 30208 5589 30245 5805
rect 30541 5589 30574 5805
rect 30208 5545 30574 5589
rect 64870 5560 64907 5856
rect 65203 5560 65252 5856
rect -3658 4731 374 4734
rect -3658 4711 454 4731
rect -3658 4255 48 4711
rect 424 4255 454 4711
rect -3658 4235 454 4255
rect -3658 4222 374 4235
rect -8372 1431 -7286 1463
rect -8372 -73 -8341 1431
rect -7317 -73 -7286 1431
rect -8372 -105 -7286 -73
rect -3650 -4316 -2690 4222
rect 13680 39 14236 61
rect 13680 35 13726 39
rect 14190 35 14236 39
rect 13680 -181 13690 35
rect 14226 -181 14236 35
rect 13680 -185 13726 -181
rect 14190 -185 14236 -181
rect 13680 -207 14236 -185
rect -3650 -4319 422 -4316
rect -3650 -4332 450 -4319
rect -3650 -4778 47 -4332
rect -8416 -5489 -7276 -5473
rect -8416 -6985 -8394 -5489
rect -7298 -5718 -7276 -5489
rect -3650 -5718 -2690 -4778
rect 20 -4788 47 -4778
rect 423 -4788 450 -4332
rect 20 -4801 450 -4788
rect 30208 -5575 30564 5545
rect 34714 4721 35132 4739
rect 31731 4710 35132 4721
rect 31731 4254 34735 4710
rect 35111 4254 35132 4710
rect 31731 4235 35132 4254
rect 31731 -4365 32061 4235
rect 34714 4225 35132 4235
rect 32542 1920 33002 1957
rect 32542 1456 32580 1920
rect 32964 1456 33002 1920
rect 32542 1419 33002 1456
rect 48466 -34 48980 -21
rect 48466 -258 48491 -34
rect 48955 -258 48980 -34
rect 48466 -271 48980 -258
rect 32560 -1506 33020 -1469
rect 32560 -1970 32598 -1506
rect 32982 -1970 33020 -1506
rect 32560 -2007 33020 -1970
rect 34726 -4321 35046 -4297
rect 34726 -4365 34738 -4321
rect 31731 -4773 34738 -4365
rect -7298 -6760 -2690 -5718
rect 30198 -5590 30578 -5575
rect 30198 -5886 30240 -5590
rect 30536 -5886 30578 -5590
rect 30198 -5901 30578 -5886
rect -7298 -6985 -7276 -6760
rect -8416 -7001 -7276 -6985
rect -3650 -14196 -2690 -6760
rect 30790 -7713 31208 -7702
rect 72 -7749 442 -7723
rect 72 -8213 105 -7749
rect 409 -8213 442 -7749
rect 72 -8239 442 -8213
rect 30790 -8417 30807 -7713
rect 31191 -7836 31208 -7713
rect 31731 -7836 32061 -4773
rect 34726 -4777 34738 -4773
rect 35034 -4777 35046 -4321
rect 34726 -4801 35046 -4777
rect 64870 -5579 65252 5560
rect 68966 4722 69424 4743
rect 68966 4698 69007 4722
rect 66018 4322 69007 4698
rect 66018 -4380 66394 4322
rect 68966 4266 69007 4322
rect 69383 4266 69424 4722
rect 68966 4245 69424 4266
rect 67036 1889 67506 1923
rect 67036 1505 67079 1889
rect 67463 1505 67506 1889
rect 67036 1471 67506 1505
rect 68976 -1502 69414 -1491
rect 68976 -1966 69003 -1502
rect 69387 -1966 69414 -1502
rect 68976 -1977 69414 -1966
rect 68976 -4312 69434 -4291
rect 68976 -4380 69017 -4312
rect 66018 -4756 69017 -4380
rect 64860 -5616 65262 -5579
rect 64860 -5992 64873 -5616
rect 65249 -5992 65262 -5616
rect 64860 -6029 65262 -5992
rect 31191 -8270 32061 -7836
rect 34730 -7767 35136 -7753
rect 34730 -8231 34741 -7767
rect 35125 -8231 35136 -7767
rect 66018 -7824 66394 -4756
rect 68976 -4768 69017 -4756
rect 69393 -4768 69434 -4312
rect 68976 -4789 69434 -4768
rect 65498 -7832 66394 -7824
rect 34730 -8245 35136 -8231
rect 65488 -7833 66394 -7832
rect 31191 -8417 31208 -8270
rect 30790 -8428 31208 -8417
rect -32 -10755 354 -10749
rect -32 -10791 13 -10755
rect 309 -10791 354 -10755
rect -32 -11175 9 -10791
rect 313 -11175 354 -10791
rect -32 -11211 13 -11175
rect 309 -11211 354 -11175
rect -32 -11217 354 -11211
rect -58 -14196 304 -14175
rect -3650 -14203 330 -14196
rect -3650 -14659 -25 -14203
rect 271 -14659 330 -14203
rect 31731 -14211 32061 -8270
rect 65488 -8297 65512 -7833
rect 65816 -8297 66394 -7833
rect 66982 -7751 67528 -7719
rect 66982 -8215 67023 -7751
rect 67487 -8215 67528 -7751
rect 66982 -8247 67528 -8215
rect 65488 -8298 66394 -8297
rect 34642 -10780 35056 -10759
rect 34642 -11244 34657 -10780
rect 35041 -11244 35056 -10780
rect 34642 -11265 35056 -11244
rect 34632 -14204 35036 -14187
rect 34632 -14211 34646 -14204
rect 31731 -14647 34646 -14211
rect -3650 -14682 330 -14659
rect 34632 -14660 34646 -14647
rect 35022 -14660 35036 -14204
rect 34632 -14677 35036 -14660
rect -3650 -14888 -2690 -14682
rect -58 -14687 304 -14682
rect 34598 -17018 35056 -16993
rect 34598 -17482 34635 -17018
rect 35019 -17482 35056 -17018
rect 34598 -17507 35056 -17482
rect 48484 -18629 48954 -18607
rect 13664 -18731 14260 -18691
rect 13664 -18875 13690 -18731
rect 14234 -18875 14260 -18731
rect 48484 -18853 48527 -18629
rect 48911 -18853 48954 -18629
rect 48484 -18875 48954 -18853
rect 13664 -18915 14260 -18875
<< via3 >>
rect 57 8162 441 8166
rect 57 7706 61 8162
rect 61 7706 437 8162
rect 437 7706 441 8162
rect 57 7702 441 7706
rect 34628 7661 34632 8285
rect 34632 7661 35168 8285
rect 35168 7661 35172 8285
rect 68987 8274 69371 8278
rect 68987 7738 68991 8274
rect 68991 7738 69367 8274
rect 69367 7738 69371 8274
rect 68987 7734 69371 7738
rect -8341 1427 -7317 1431
rect -8341 -69 -8337 1427
rect -8337 -69 -7321 1427
rect -7321 -69 -7317 1427
rect -8341 -73 -7317 -69
rect 13726 35 14190 39
rect 13726 -181 14190 35
rect 13726 -185 14190 -181
rect 32580 1916 32964 1920
rect 32580 1460 32584 1916
rect 32584 1460 32960 1916
rect 32960 1460 32964 1916
rect 32580 1456 32964 1460
rect 48491 -38 48955 -34
rect 48491 -254 48495 -38
rect 48495 -254 48951 -38
rect 48951 -254 48955 -38
rect 48491 -258 48955 -254
rect 32598 -1510 32982 -1506
rect 32598 -1966 32602 -1510
rect 32602 -1966 32978 -1510
rect 32978 -1966 32982 -1510
rect 32598 -1970 32982 -1966
rect 105 -7753 409 -7749
rect 105 -8209 109 -7753
rect 109 -8209 405 -7753
rect 405 -8209 409 -7753
rect 105 -8213 409 -8209
rect 30807 -8417 31191 -7713
rect 67079 1885 67463 1889
rect 67079 1509 67083 1885
rect 67083 1509 67459 1885
rect 67459 1509 67463 1885
rect 67079 1505 67463 1509
rect 69003 -1506 69387 -1502
rect 69003 -1962 69007 -1506
rect 69007 -1962 69383 -1506
rect 69383 -1962 69387 -1506
rect 69003 -1966 69387 -1962
rect 34741 -7771 35125 -7767
rect 34741 -8227 34745 -7771
rect 34745 -8227 35121 -7771
rect 35121 -8227 35125 -7771
rect 34741 -8231 35125 -8227
rect 9 -11175 13 -10791
rect 13 -11175 309 -10791
rect 309 -11175 313 -10791
rect 65512 -8297 65816 -7833
rect 67023 -7755 67487 -7751
rect 67023 -8211 67027 -7755
rect 67027 -8211 67483 -7755
rect 67483 -8211 67487 -7755
rect 67023 -8215 67487 -8211
rect 34657 -10784 35041 -10780
rect 34657 -11240 34661 -10784
rect 34661 -11240 35037 -10784
rect 35037 -11240 35041 -10784
rect 34657 -11244 35041 -11240
rect 34635 -17022 35019 -17018
rect 34635 -17478 34639 -17022
rect 34639 -17478 35015 -17022
rect 35015 -17478 35019 -17022
rect 34635 -17482 35019 -17478
rect 13690 -18735 14234 -18731
rect 13690 -18871 13694 -18735
rect 13694 -18871 14230 -18735
rect 14230 -18871 14234 -18735
rect 13690 -18875 14234 -18871
rect 48527 -18633 48911 -18629
rect 48527 -18849 48531 -18633
rect 48531 -18849 48907 -18633
rect 48907 -18849 48911 -18633
rect 48527 -18853 48911 -18849
<< metal4 >>
rect 34617 8285 35183 8323
rect 34617 8232 34628 8285
rect 43 8168 455 8191
rect -1944 8166 461 8168
rect -1944 8139 57 8166
rect -1945 7706 57 8139
rect -8363 1431 -7295 1459
rect -8363 -73 -8341 1431
rect -7317 1170 -7295 1431
rect -1945 1170 -959 7706
rect 43 7702 57 7706
rect 441 7706 461 8166
rect 30744 7770 34628 8232
rect 441 7702 455 7706
rect 43 7677 455 7702
rect 32562 1953 33002 1966
rect 32551 1920 33002 1953
rect 32551 1456 32580 1920
rect 32964 1456 33002 1920
rect 32551 1423 33002 1456
rect -7317 120 -959 1170
rect -7317 106 -6654 120
rect -7317 -73 -7295 106
rect -8363 -101 -7295 -73
rect -1945 -1494 -959 120
rect 13689 45 14227 57
rect 13689 39 13840 45
rect 14076 39 14227 45
rect 13689 -185 13726 39
rect 14190 -185 14227 39
rect 13689 -191 13840 -185
rect 14076 -191 14227 -185
rect 13689 -203 14227 -191
rect 32562 -1473 33002 1423
rect -1945 -1974 -956 -1494
rect 32562 -1506 33011 -1473
rect 32562 -1970 32598 -1506
rect 32982 -1970 33011 -1506
rect -1945 -7746 -959 -1974
rect 32562 -2003 33011 -1970
rect 30799 -7713 31199 -7701
rect 81 -7746 433 -7727
rect -1945 -7749 433 -7746
rect -1945 -8213 105 -7749
rect 409 -8213 433 -7749
rect -1945 -8235 433 -8213
rect -1945 -8252 424 -8235
rect -1945 -10754 -959 -8252
rect 30799 -8417 30807 -7713
rect 31191 -8417 31199 -7713
rect 30799 -8429 31199 -8417
rect 32562 -10702 33002 -2003
rect -23 -10754 345 -10753
rect -1945 -10791 368 -10754
rect -1945 -11175 9 -10791
rect 313 -11175 368 -10791
rect 30724 -11170 33002 -10702
rect -1945 -11244 368 -11175
rect -1945 -11349 -959 -11244
rect 32562 -17048 33002 -11170
rect 33501 -7779 33963 7770
rect 34617 7661 34628 7770
rect 35172 7661 35183 8285
rect 68961 8278 69397 8283
rect 68961 8230 68987 8278
rect 65430 7768 68987 8230
rect 34617 7623 35183 7661
rect 67039 1889 67501 2069
rect 67039 1505 67079 1889
rect 67463 1505 67501 1889
rect 48472 -20 48974 -16
rect 48472 -34 48605 -20
rect 48841 -34 48974 -20
rect 48472 -258 48491 -34
rect 48955 -258 48974 -34
rect 48472 -260 48974 -258
rect 48475 -267 48971 -260
rect 67039 -7723 67501 1505
rect 68099 -1481 68561 7768
rect 68961 7734 68987 7768
rect 69371 7734 69397 8278
rect 68961 7729 69397 7734
rect 99684 2343 100146 8234
rect 101138 2343 102002 3218
rect 99684 1881 102002 2343
rect 101138 1068 102002 1881
rect 68099 -1495 69367 -1481
rect 68099 -1502 69405 -1495
rect 68099 -1943 69003 -1502
rect 68985 -1966 69003 -1943
rect 69387 -1966 69405 -1502
rect 68985 -1973 69405 -1966
rect 66991 -7751 67519 -7723
rect 34739 -7767 35127 -7757
rect 34739 -7779 34741 -7767
rect 33501 -8231 34741 -7779
rect 35125 -8231 35127 -7767
rect 33501 -8241 35127 -8231
rect 65497 -7833 65831 -7831
rect 33501 -10785 33963 -8241
rect 65497 -8297 65512 -7833
rect 65816 -8297 65831 -7833
rect 66991 -8215 67023 -7751
rect 67487 -8215 67519 -7751
rect 101154 -7811 102018 -7008
rect 66991 -8243 67519 -8215
rect 65497 -8299 65831 -8297
rect 67039 -10696 67501 -8243
rect 99678 -8273 102018 -7811
rect 101154 -9158 102018 -8273
rect 34651 -10780 35047 -10763
rect 34651 -10785 34657 -10780
rect 33501 -11244 34657 -10785
rect 35041 -11244 35047 -10780
rect 65334 -11158 67663 -10696
rect 33501 -11247 35047 -11244
rect 34651 -11261 35047 -11247
rect 34607 -17018 35047 -16997
rect 34607 -17048 34635 -17018
rect 32562 -17482 34635 -17048
rect 35019 -17482 35047 -17018
rect 32562 -17488 35047 -17482
rect 34607 -17503 35047 -17488
rect 13684 -18601 14224 -18550
rect 13684 -18695 13836 -18601
rect 13673 -18731 13836 -18695
rect 14072 -18695 14224 -18601
rect 48493 -18623 48945 -18611
rect 48493 -18629 48601 -18623
rect 48837 -18629 48945 -18623
rect 14072 -18731 14251 -18695
rect 13673 -18875 13690 -18731
rect 14234 -18875 14251 -18731
rect 48493 -18853 48527 -18629
rect 48911 -18853 48945 -18629
rect 48493 -18859 48601 -18853
rect 48837 -18859 48945 -18853
rect 48493 -18871 48945 -18859
rect 13673 -18911 14251 -18875
<< via4 >>
rect 13840 39 14076 45
rect 13840 -185 14076 39
rect 13840 -191 14076 -185
rect 48605 -34 48841 -20
rect 48605 -256 48841 -34
rect 13836 -18731 14072 -18601
rect 48601 -18629 48837 -18623
rect 13836 -18837 14072 -18731
rect 48601 -18853 48837 -18629
rect 48601 -18859 48837 -18853
<< metal5 >>
rect 13662 45 14254 100
rect 13662 -191 13840 45
rect 14076 -191 14254 45
rect 13662 -382 14254 -191
rect 48444 -20 49002 10
rect 48444 -256 48605 -20
rect 48841 -256 49002 -20
rect 48444 -362 49002 -256
rect 13674 -18526 14244 -382
rect 13660 -18601 14248 -18526
rect 13660 -18837 13836 -18601
rect 14072 -18837 14248 -18601
rect 48452 -18623 48996 -362
rect 48452 -18672 48601 -18623
rect 13660 -18912 14248 -18837
rect 48454 -18859 48601 -18672
rect 48837 -18672 48996 -18623
rect 48837 -18859 48994 -18672
rect 48454 -18904 48994 -18859
use analog_neuron_3input_re  analog_neuron_3input_re_1
timestamp 1627926120
transform 1 0 460 0 1 -12660
box -548 -6266 30658 3151
use sky130_fd_pr__res_xhigh_po_0p35_95A2JL  sky130_fd_pr__res_xhigh_po_0p35_95A2JL_0
timestamp 1627926120
transform 0 1 17195 -1 0 -14333
box -35 -1325 35 1325
use sky130_fd_pr__res_xhigh_po_0p35_S33692  sky130_fd_pr__res_xhigh_po_0p35_S33692_0
timestamp 1627926120
transform 0 1 17065 -1 0 -15551
box -35 -531 35 531
use sky130_fd_pr__res_high_po_0p35_AXF3YZ  sky130_fd_pr__res_high_po_0p35_AXF3YZ_0
timestamp 1627926120
transform 0 1 17152 -1 0 -16853
box -35 -694 35 694
use analog_neuron_3input_re  analog_neuron_3input_re_3
timestamp 1627926120
transform 1 0 35146 0 1 -12662
box -548 -6266 30658 3151
use sky130_fd_pr__res_high_po_0p35_8YJL8A  sky130_fd_pr__res_high_po_0p35_8YJL8A_0
timestamp 1627926120
transform 0 1 51781 -1 0 -14349
box -35 -1037 35 1037
use sky130_fd_pr__res_high_po_0p35_PMTBZG  sky130_fd_pr__res_high_po_0p35_PMTBZG_0
timestamp 1627926120
transform 0 1 51527 -1 0 -16853
box -35 -967 35 967
use analog_neuron_3input_re  analog_neuron_3input_re_0
timestamp 1627926120
transform 1 0 550 0 -1 -6309
box -548 -6266 30658 3151
use analog_neuron_3input_re  analog_neuron_3input_re_2
timestamp 1627926120
transform 1 0 35236 0 -1 -6311
box -548 -6266 30658 3151
use sky130_fd_pr__res_xhigh_po_0p35_KDN527  sky130_fd_pr__res_xhigh_po_0p35_KDN527_0
timestamp 1627926120
transform 0 1 86055 -1 0 -2135
box -35 -683 35 683
use analog_neuron_3input_re  analog_neuron_3input_re_4
timestamp 1627926120
transform 1 0 69490 0 -1 -6307
box -548 -6266 30658 3151
use sky130_fd_pr__res_xhigh_po_0p35_X3XLR2  sky130_fd_pr__res_xhigh_po_0p35_X3XLR2_0
timestamp 1627926120
transform 0 1 17241 -1 0 4579
box -35 -1267 35 1267
use analog_neuron_3input_re  analog_neuron_3input_re_5
timestamp 1627926120
transform 1 0 548 0 1 6266
box -548 -6266 30658 3151
use sky130_fd_pr__res_xhigh_po_0p35_MT7BFK  sky130_fd_pr__res_xhigh_po_0p35_MT7BFK_0
timestamp 1627926120
transform 0 1 17075 -1 0 3345
box -35 -541 35 541
use sky130_fd_pr__res_high_po_0p35_4RFVXF  sky130_fd_pr__res_high_po_0p35_4RFVXF_0
timestamp 1627926120
transform 0 1 17246 -1 0 2097
box -35 -724 35 724
use analog_neuron_3input_re  analog_neuron_3input_re_6
timestamp 1627926120
transform 1 0 35234 0 1 6264
box -548 -6266 30658 3151
use sky130_fd_pr__res_xhigh_po_0p35_T8PEF7  sky130_fd_pr__res_xhigh_po_0p35_T8PEF7_0
timestamp 1627926120
transform 0 1 51782 -1 0 4586
box -35 -815 35 815
use sky130_fd_pr__res_xhigh_po_0p35_RG46CN  sky130_fd_pr__res_xhigh_po_0p35_RG46CN_0
timestamp 1627926120
transform 0 1 51881 -1 0 2099
box -35 -775 35 775
use analog_neuron_3input_re  analog_neuron_3input_re_7
timestamp 1627926120
transform 1 0 69488 0 1 6268
box -548 -6266 30658 3151
use sky130_fd_pr__res_xhigh_po_0p35_M9RFTX  sky130_fd_pr__res_xhigh_po_0p35_M9RFTX_0
timestamp 1627926120
transform 0 1 86138 -1 0 4563
box -35 -1070 35 1070
use sky130_fd_pr__res_xhigh_po_0p35_7NH2RC  sky130_fd_pr__res_xhigh_po_0p35_7NH2RC_0
timestamp 1627926120
transform 0 1 86152 -1 0 2063
box -35 -712 35 712
<< labels >>
rlabel metal4 s 101282 -9094 101942 -7102 4 Out2
port 1 nsew
rlabel metal4 s 101208 1120 101868 3112 4 Out1
port 2 nsew
rlabel metal2 s -8490 -382 -7204 1836 4 In1
port 3 nsew
rlabel metal2 s -8528 -7322 -7242 -5104 4 In2
port 4 nsew
rlabel metal2 s -8472 -13574 -7186 -11356 4 In3
port 5 nsew
rlabel metal2 s 1472 9288 99492 9404 4 VDD
port 6 nsew
rlabel metal2 s 4408 -9582 36564 -9412 4 VDD
port 6 nsew
rlabel metal2 s 38920 -9594 99424 -9412 4 VDD
port 6 nsew
rlabel metal2 s 2048 -18912 63536 -18810 4 GND
port 7 nsew
rlabel metal2 s 21232 -132 54090 64 4 GND
port 7 nsew
rlabel metal2 s 55578 -140 88294 60 4 GND
port 7 nsew
rlabel metal2 s 89822 -154 97866 90 4 GND
port 7 nsew
rlabel metal2 s 2040 -138 19166 102 4 GND
port 7 nsew
<< end >>
