magic
tech sky130A
magscale 1 2
timestamp 1628283727
<< xpolycontact >>
rect -69 96 69 528
rect -69 -528 69 -96
<< ppolyres >>
rect -69 -96 69 96
<< viali >>
rect -53 113 53 510
rect -53 -510 53 -113
<< metal1 >>
rect -59 510 59 522
rect -59 113 -53 510
rect 53 113 59 510
rect -59 101 59 113
rect -59 -113 59 -101
rect -59 -510 -53 -113
rect 53 -510 59 -113
rect -59 -522 59 -510
<< res0p69 >>
rect -71 -98 71 98
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p69
string parameters w 0.690 l .96 m 1 nx 1 wmin 0.690 lmin 0.50 rho 319.8 val 500.556 dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
