magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 109 35 541
rect -35 -541 35 -109
<< xpolyres >>
rect -35 -109 35 109
<< viali >>
rect -17 487 17 521
rect -17 415 17 449
rect -17 343 17 377
rect -17 271 17 305
rect -17 199 17 233
rect -17 127 17 161
rect -17 -162 17 -128
rect -17 -234 17 -200
rect -17 -306 17 -272
rect -17 -378 17 -344
rect -17 -450 17 -416
rect -17 -522 17 -488
<< metal1 >>
rect -25 521 25 535
rect -25 487 -17 521
rect 17 487 25 521
rect -25 449 25 487
rect -25 415 -17 449
rect 17 415 25 449
rect -25 377 25 415
rect -25 343 -17 377
rect 17 343 25 377
rect -25 305 25 343
rect -25 271 -17 305
rect 17 271 25 305
rect -25 233 25 271
rect -25 199 -17 233
rect 17 199 25 233
rect -25 161 25 199
rect -25 127 -17 161
rect 17 127 25 161
rect -25 114 25 127
rect -25 -128 25 -114
rect -25 -162 -17 -128
rect 17 -162 25 -128
rect -25 -200 25 -162
rect -25 -234 -17 -200
rect 17 -234 25 -200
rect -25 -272 25 -234
rect -25 -306 -17 -272
rect 17 -306 25 -272
rect -25 -344 25 -306
rect -25 -378 -17 -344
rect 17 -378 25 -344
rect -25 -416 25 -378
rect -25 -450 -17 -416
rect 17 -450 25 -416
rect -25 -488 25 -450
rect -25 -522 -17 -488
rect 17 -522 25 -488
rect -25 -535 25 -522
<< end >>
