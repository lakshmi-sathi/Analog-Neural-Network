magic
tech sky130A
magscale 1 2
timestamp 1627921586
<< xpolycontact >>
rect -35 109 35 541
rect -35 -541 35 -109
<< xpolyres >>
rect -35 -109 35 109
<< viali >>
rect -19 126 19 523
rect -19 -523 19 -126
<< metal1 >>
rect -25 523 25 535
rect -25 126 -19 523
rect 19 126 25 523
rect -25 114 25 126
rect -25 -126 25 -114
rect -25 -523 -19 -126
rect 19 -523 25 -126
rect -25 -535 25 -523
<< res0p35 >>
rect -37 -111 37 111
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 1.09 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 6.914k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
