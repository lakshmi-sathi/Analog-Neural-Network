magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< nwell >>
rect 518 1248 582 1268
rect 710 1248 774 1264
rect 902 1248 966 1266
rect 518 1222 612 1248
rect 518 1208 596 1222
rect 710 1218 804 1248
rect 902 1220 996 1248
rect 710 1208 786 1218
rect 902 1208 980 1220
rect 518 1118 582 1208
rect 710 1114 774 1208
rect 902 1116 966 1208
rect 1094 1120 1158 1270
rect 612 332 684 566
rect 604 292 684 332
rect 678 148 708 158
rect 870 148 900 158
rect 564 96 1030 148
rect 1062 142 1092 158
<< poly >>
rect 1062 105 1092 151
rect 1009 101 1092 105
rect 997 75 1092 101
<< locali >>
rect 478 1388 1194 1408
rect 478 1354 498 1388
rect 532 1354 570 1388
rect 604 1354 642 1388
rect 676 1354 714 1388
rect 748 1354 786 1388
rect 820 1354 858 1388
rect 892 1354 930 1388
rect 964 1354 1002 1388
rect 1036 1354 1074 1388
rect 1108 1354 1146 1388
rect 1180 1354 1194 1388
rect 478 1336 1194 1354
rect -38 -46 46 10
<< viali >>
rect 498 1354 532 1388
rect 570 1354 604 1388
rect 642 1354 676 1388
rect 714 1354 748 1388
rect 786 1354 820 1388
rect 858 1354 892 1388
rect 930 1354 964 1388
rect 1002 1354 1036 1388
rect 1074 1354 1108 1388
rect 1146 1354 1180 1388
<< metal1 >>
rect 482 1397 1188 1404
rect 482 1388 555 1397
rect 482 1354 498 1388
rect 532 1354 555 1388
rect 482 1345 555 1354
rect 607 1345 619 1397
rect 671 1388 683 1397
rect 735 1388 747 1397
rect 799 1388 811 1397
rect 863 1388 875 1397
rect 927 1388 939 1397
rect 991 1388 1003 1397
rect 676 1354 683 1388
rect 927 1354 930 1388
rect 991 1354 1002 1388
rect 671 1345 683 1354
rect 735 1345 747 1354
rect 799 1345 811 1354
rect 863 1345 875 1354
rect 927 1345 939 1354
rect 991 1345 1003 1354
rect 1055 1345 1067 1397
rect 1119 1388 1188 1397
rect 1119 1354 1146 1388
rect 1180 1354 1188 1388
rect 1119 1345 1188 1354
rect 482 1336 1188 1345
rect 128 1222 190 1276
rect 656 1202 1120 1250
rect 68 1158 142 1184
rect 68 1106 76 1158
rect 128 1106 142 1158
rect 68 1094 142 1106
rect 68 1042 76 1094
rect 128 1042 142 1094
rect 68 1030 142 1042
rect 68 978 76 1030
rect 128 978 142 1030
rect 68 966 142 978
rect 68 914 76 966
rect 128 914 142 966
rect 68 902 142 914
rect 68 850 76 902
rect 128 850 142 902
rect 68 838 142 850
rect 68 786 76 838
rect 128 786 142 838
rect 518 1141 582 1174
rect 518 1089 524 1141
rect 576 1089 582 1141
rect 518 1077 582 1089
rect 518 1025 524 1077
rect 576 1025 582 1077
rect 518 1013 582 1025
rect 518 961 524 1013
rect 576 961 582 1013
rect 518 949 582 961
rect 518 897 524 949
rect 576 897 582 949
rect 518 885 582 897
rect 518 833 524 885
rect 576 833 582 885
rect 518 808 582 833
rect 710 1151 774 1174
rect 710 1099 716 1151
rect 768 1099 774 1151
rect 710 1087 774 1099
rect 710 1035 716 1087
rect 768 1035 774 1087
rect 710 1023 774 1035
rect 710 971 716 1023
rect 768 971 774 1023
rect 710 959 774 971
rect 710 907 716 959
rect 768 907 774 959
rect 710 895 774 907
rect 710 843 716 895
rect 768 843 774 895
rect 710 828 774 843
rect 902 1154 966 1174
rect 902 1102 908 1154
rect 960 1102 966 1154
rect 902 1090 966 1102
rect 902 1038 908 1090
rect 960 1038 966 1090
rect 902 1026 966 1038
rect 902 974 908 1026
rect 960 974 966 1026
rect 902 962 966 974
rect 902 910 908 962
rect 960 910 966 962
rect 902 898 966 910
rect 902 846 908 898
rect 960 846 966 898
rect 902 834 966 846
rect 1094 1140 1158 1174
rect 1094 1088 1100 1140
rect 1152 1088 1158 1140
rect 1094 1076 1158 1088
rect 1094 1024 1100 1076
rect 1152 1024 1158 1076
rect 1094 1012 1158 1024
rect 1094 960 1100 1012
rect 1152 960 1158 1012
rect 1094 948 1158 960
rect 1094 896 1100 948
rect 1152 896 1158 948
rect 1094 884 1158 896
rect 1094 832 1100 884
rect 1152 832 1158 884
rect 1094 806 1158 832
rect 68 768 142 786
rect 174 546 240 556
rect 174 494 180 546
rect 232 494 240 546
rect 174 482 240 494
rect 174 430 180 482
rect 232 430 240 482
rect 174 418 240 430
rect 174 366 180 418
rect 232 366 240 418
rect 174 354 240 366
rect 174 302 180 354
rect 232 302 240 354
rect 174 290 240 302
rect 174 238 180 290
rect 232 238 240 290
rect 174 226 240 238
rect 174 174 180 226
rect 232 174 240 226
rect 174 158 240 174
rect 614 509 680 540
rect 614 457 620 509
rect 672 457 680 509
rect 614 445 680 457
rect 614 393 620 445
rect 672 393 680 445
rect 614 381 680 393
rect 614 329 620 381
rect 672 329 680 381
rect 614 317 680 329
rect 614 265 620 317
rect 672 265 680 317
rect 614 253 680 265
rect 614 201 620 253
rect 672 201 680 253
rect 614 164 680 201
rect 806 509 872 540
rect 806 457 812 509
rect 864 457 872 509
rect 806 445 872 457
rect 806 393 812 445
rect 864 393 872 445
rect 806 381 872 393
rect 806 329 812 381
rect 864 329 872 381
rect 806 317 872 329
rect 806 265 812 317
rect 864 265 872 317
rect 806 253 872 265
rect 806 201 812 253
rect 864 201 872 253
rect 806 164 872 201
rect 998 508 1064 538
rect 998 456 1004 508
rect 1056 456 1064 508
rect 998 444 1064 456
rect 998 392 1004 444
rect 1056 392 1064 444
rect 998 380 1064 392
rect 998 328 1004 380
rect 1056 328 1064 380
rect 998 316 1064 328
rect 998 264 1004 316
rect 1056 264 1064 316
rect 998 252 1064 264
rect 998 200 1004 252
rect 1056 200 1064 252
rect 998 164 1064 200
rect 564 120 1030 122
rect -102 32 1030 120
<< via1 >>
rect 555 1388 607 1397
rect 555 1354 570 1388
rect 570 1354 604 1388
rect 604 1354 607 1388
rect 555 1345 607 1354
rect 619 1388 671 1397
rect 683 1388 735 1397
rect 747 1388 799 1397
rect 811 1388 863 1397
rect 875 1388 927 1397
rect 939 1388 991 1397
rect 1003 1388 1055 1397
rect 619 1354 642 1388
rect 642 1354 671 1388
rect 683 1354 714 1388
rect 714 1354 735 1388
rect 747 1354 748 1388
rect 748 1354 786 1388
rect 786 1354 799 1388
rect 811 1354 820 1388
rect 820 1354 858 1388
rect 858 1354 863 1388
rect 875 1354 892 1388
rect 892 1354 927 1388
rect 939 1354 964 1388
rect 964 1354 991 1388
rect 1003 1354 1036 1388
rect 1036 1354 1055 1388
rect 619 1345 671 1354
rect 683 1345 735 1354
rect 747 1345 799 1354
rect 811 1345 863 1354
rect 875 1345 927 1354
rect 939 1345 991 1354
rect 1003 1345 1055 1354
rect 1067 1388 1119 1397
rect 1067 1354 1074 1388
rect 1074 1354 1108 1388
rect 1108 1354 1119 1388
rect 1067 1345 1119 1354
rect 76 1106 128 1158
rect 76 1042 128 1094
rect 76 978 128 1030
rect 76 914 128 966
rect 76 850 128 902
rect 76 786 128 838
rect 524 1089 576 1141
rect 524 1025 576 1077
rect 524 961 576 1013
rect 524 897 576 949
rect 524 833 576 885
rect 716 1099 768 1151
rect 716 1035 768 1087
rect 716 971 768 1023
rect 716 907 768 959
rect 716 843 768 895
rect 908 1102 960 1154
rect 908 1038 960 1090
rect 908 974 960 1026
rect 908 910 960 962
rect 908 846 960 898
rect 1100 1088 1152 1140
rect 1100 1024 1152 1076
rect 1100 960 1152 1012
rect 1100 896 1152 948
rect 1100 832 1152 884
rect 180 494 232 546
rect 180 430 232 482
rect 180 366 232 418
rect 180 302 232 354
rect 180 238 232 290
rect 180 174 232 226
rect 620 457 672 509
rect 620 393 672 445
rect 620 329 672 381
rect 620 265 672 317
rect 620 201 672 253
rect 812 457 864 509
rect 812 393 864 445
rect 812 329 864 381
rect 812 265 864 317
rect 812 201 864 253
rect 1004 456 1056 508
rect 1004 392 1056 444
rect 1004 328 1056 380
rect 1004 264 1056 316
rect 1004 200 1056 252
<< metal2 >>
rect -50 1426 1308 1530
rect 518 1397 1158 1426
rect 518 1345 555 1397
rect 607 1345 619 1397
rect 671 1345 683 1397
rect 735 1345 747 1397
rect 799 1345 811 1397
rect 863 1345 875 1397
rect 927 1345 939 1397
rect 991 1345 1003 1397
rect 1055 1345 1067 1397
rect 1119 1345 1158 1397
rect 518 1262 1158 1345
rect 68 1158 142 1184
rect 68 1106 76 1158
rect 128 1106 142 1158
rect 68 1094 142 1106
rect 68 1042 76 1094
rect 128 1042 142 1094
rect 68 1030 142 1042
rect 68 978 76 1030
rect 128 978 142 1030
rect 68 966 142 978
rect 68 914 76 966
rect 128 914 142 966
rect 68 902 142 914
rect 68 859 76 902
rect -25 850 76 859
rect 128 850 142 902
rect -25 838 142 850
rect -25 786 76 838
rect 128 786 142 838
rect 518 1141 582 1262
rect 518 1089 524 1141
rect 576 1089 582 1141
rect 518 1077 582 1089
rect 518 1025 524 1077
rect 576 1025 582 1077
rect 518 1013 582 1025
rect 518 961 524 1013
rect 576 961 582 1013
rect 518 949 582 961
rect 518 897 524 949
rect 576 897 582 949
rect 518 885 582 897
rect 518 833 524 885
rect 576 833 582 885
rect 518 808 582 833
rect 710 1151 774 1262
rect 710 1099 716 1151
rect 768 1099 774 1151
rect 710 1087 774 1099
rect 710 1035 716 1087
rect 768 1035 774 1087
rect 710 1023 774 1035
rect 710 971 716 1023
rect 768 971 774 1023
rect 710 959 774 971
rect 710 907 716 959
rect 768 907 774 959
rect 710 895 774 907
rect 710 843 716 895
rect 768 843 774 895
rect 710 828 774 843
rect 902 1154 966 1262
rect 902 1102 908 1154
rect 960 1102 966 1154
rect 902 1090 966 1102
rect 902 1038 908 1090
rect 960 1038 966 1090
rect 902 1026 966 1038
rect 902 974 908 1026
rect 960 974 966 1026
rect 902 962 966 974
rect 902 910 908 962
rect 960 910 966 962
rect 902 898 966 910
rect 902 846 908 898
rect 960 846 966 898
rect 902 834 966 846
rect 1094 1140 1158 1262
rect 1094 1088 1100 1140
rect 1152 1088 1158 1140
rect 1094 1076 1158 1088
rect 1094 1024 1100 1076
rect 1152 1024 1158 1076
rect 1094 1012 1158 1024
rect 1094 960 1100 1012
rect 1152 960 1158 1012
rect 1094 948 1158 960
rect 1094 896 1100 948
rect 1152 896 1158 948
rect 1094 884 1158 896
rect 1094 832 1100 884
rect 1152 832 1158 884
rect 1094 806 1158 832
rect -25 768 142 786
rect -25 763 141 768
rect -25 -66 37 763
rect 174 552 240 566
rect 174 494 180 552
rect 236 496 240 552
rect 614 540 680 550
rect 232 494 240 496
rect 174 482 240 494
rect 174 238 180 482
rect 232 472 240 482
rect 236 416 240 472
rect 232 392 240 416
rect 236 336 240 392
rect 232 312 240 336
rect 236 256 240 312
rect 232 238 240 256
rect 174 232 240 238
rect 174 174 180 232
rect 236 176 240 232
rect 232 174 240 176
rect 174 158 240 174
rect 612 509 680 540
rect 612 505 620 509
rect 672 505 680 509
rect 612 449 618 505
rect 674 449 680 505
rect 612 445 680 449
rect 612 425 620 445
rect 672 425 680 445
rect 612 369 618 425
rect 674 369 680 425
rect 612 345 620 369
rect 672 345 680 369
rect 612 289 618 345
rect 674 289 680 345
rect 612 265 620 289
rect 672 265 680 289
rect 612 209 618 265
rect 674 209 680 265
rect 612 201 620 209
rect 672 201 680 209
rect 612 160 680 201
rect 804 509 872 550
rect 804 505 812 509
rect 864 505 872 509
rect 804 449 810 505
rect 866 449 872 505
rect 804 445 872 449
rect 804 425 812 445
rect 864 425 872 445
rect 804 369 810 425
rect 866 369 872 425
rect 804 345 812 369
rect 864 345 872 369
rect 804 289 810 345
rect 866 289 872 345
rect 804 265 812 289
rect 864 265 872 289
rect 804 209 810 265
rect 866 209 872 265
rect 804 201 812 209
rect 864 201 872 209
rect 804 160 872 201
rect 996 508 1064 550
rect 996 504 1004 508
rect 1056 504 1064 508
rect 996 448 1002 504
rect 1058 448 1064 504
rect 996 444 1064 448
rect 996 424 1004 444
rect 1056 424 1064 444
rect 996 368 1002 424
rect 1058 368 1064 424
rect 996 344 1004 368
rect 1056 344 1064 368
rect 996 288 1002 344
rect 1058 288 1064 344
rect 996 264 1004 288
rect 1056 264 1064 288
rect 996 208 1002 264
rect 1058 208 1064 264
rect 996 200 1004 208
rect 1056 200 1064 208
rect 996 160 1064 200
rect -58 -170 1300 -66
<< via2 >>
rect 180 546 236 552
rect 180 496 232 546
rect 232 496 236 546
rect 180 430 232 472
rect 232 430 236 472
rect 180 418 236 430
rect 180 416 232 418
rect 232 416 236 418
rect 180 366 232 392
rect 232 366 236 392
rect 180 354 236 366
rect 180 336 232 354
rect 232 336 236 354
rect 180 302 232 312
rect 232 302 236 312
rect 180 290 236 302
rect 180 256 232 290
rect 232 256 236 290
rect 180 226 236 232
rect 180 176 232 226
rect 232 176 236 226
rect 618 457 620 505
rect 620 457 672 505
rect 672 457 674 505
rect 618 449 674 457
rect 618 393 620 425
rect 620 393 672 425
rect 672 393 674 425
rect 618 381 674 393
rect 618 369 620 381
rect 620 369 672 381
rect 672 369 674 381
rect 618 329 620 345
rect 620 329 672 345
rect 672 329 674 345
rect 618 317 674 329
rect 618 289 620 317
rect 620 289 672 317
rect 672 289 674 317
rect 618 253 674 265
rect 618 209 620 253
rect 620 209 672 253
rect 672 209 674 253
rect 810 457 812 505
rect 812 457 864 505
rect 864 457 866 505
rect 810 449 866 457
rect 810 393 812 425
rect 812 393 864 425
rect 864 393 866 425
rect 810 381 866 393
rect 810 369 812 381
rect 812 369 864 381
rect 864 369 866 381
rect 810 329 812 345
rect 812 329 864 345
rect 864 329 866 345
rect 810 317 866 329
rect 810 289 812 317
rect 812 289 864 317
rect 864 289 866 317
rect 810 253 866 265
rect 810 209 812 253
rect 812 209 864 253
rect 864 209 866 253
rect 1002 456 1004 504
rect 1004 456 1056 504
rect 1056 456 1058 504
rect 1002 448 1058 456
rect 1002 392 1004 424
rect 1004 392 1056 424
rect 1056 392 1058 424
rect 1002 380 1058 392
rect 1002 368 1004 380
rect 1004 368 1056 380
rect 1056 368 1058 380
rect 1002 328 1004 344
rect 1004 328 1056 344
rect 1056 328 1058 344
rect 1002 316 1058 328
rect 1002 288 1004 316
rect 1004 288 1056 316
rect 1056 288 1058 316
rect 1002 252 1058 264
rect 1002 208 1004 252
rect 1004 208 1056 252
rect 1056 208 1058 252
<< metal3 >>
rect 174 556 242 566
rect 172 552 250 556
rect 172 496 180 552
rect 236 496 250 552
rect 172 472 250 496
rect 172 416 180 472
rect 236 416 250 472
rect 172 392 250 416
rect 172 336 180 392
rect 236 336 250 392
rect 172 312 250 336
rect 172 304 180 312
rect 174 256 180 304
rect 236 256 250 312
rect 174 232 250 256
rect 174 176 180 232
rect 236 212 250 232
rect 612 540 682 550
rect 804 540 872 550
rect 612 505 684 540
rect 612 449 618 505
rect 674 449 684 505
rect 612 425 684 449
rect 612 369 618 425
rect 674 369 684 425
rect 612 345 684 369
rect 612 289 618 345
rect 674 306 684 345
rect 802 505 872 540
rect 996 538 1064 550
rect 802 449 810 505
rect 866 449 872 505
rect 802 425 872 449
rect 802 369 810 425
rect 866 369 872 425
rect 802 345 872 369
rect 802 306 810 345
rect 674 289 682 306
rect 612 265 682 289
rect 612 212 618 265
rect 236 209 618 212
rect 674 212 682 265
rect 804 289 810 306
rect 866 289 872 345
rect 804 265 872 289
rect 804 212 810 265
rect 674 209 810 212
rect 866 212 872 265
rect 994 504 1064 538
rect 994 448 1002 504
rect 1058 448 1064 504
rect 994 424 1064 448
rect 994 368 1002 424
rect 1058 368 1064 424
rect 994 350 1064 368
rect 994 344 1068 350
rect 994 288 1002 344
rect 1058 288 1068 344
rect 994 264 1068 288
rect 994 212 1002 264
rect 866 209 1002 212
rect 236 208 1002 209
rect 1058 212 1068 264
rect 1058 208 1308 212
rect 236 176 1308 208
rect 174 118 1308 176
rect 174 116 1292 118
use sky130_fd_pr__pfet_01v8_27F7GK  sky130_fd_pr__pfet_01v8_27F7GK_0
timestamp 1627926120
transform 1 0 837 0 1 661
box -455 -719 455 719
use sky130_fd_pr__nfet_01v8_LW2HKK  sky130_fd_pr__nfet_01v8_LW2HKK_0
timestamp 1627926120
transform 1 0 161 0 1 670
box -175 -694 175 694
<< labels >>
rlabel metal1 s -102 32 -28 120 4 in
port 1 nsew
rlabel metal2 s -44 1430 1302 1524 4 vh
port 2 nsew
rlabel metal2 s -54 -164 1294 -72 4 vl
port 3 nsew
rlabel locali s -32 -40 40 4 4 nbody
port 4 nsew
rlabel metal3 s 1208 122 1304 208 4 out
port 5 nsew
<< end >>
