magic
tech sky130A
magscale 1 2
timestamp 1627111729
<< error_p >>
rect -29 129 29 135
rect -29 95 -17 129
rect -29 89 29 95
<< nwell >>
rect -109 -182 109 148
<< pmos >>
rect -15 -120 15 48
<< pdiff >>
rect -73 36 -15 48
rect -73 -108 -61 36
rect -27 -108 -15 36
rect -73 -120 -15 -108
rect 15 36 73 48
rect 15 -108 27 36
rect 61 -108 73 36
rect 15 -120 73 -108
<< pdiffc >>
rect -61 -108 -27 36
rect 27 -108 61 36
<< poly >>
rect -33 129 33 145
rect -33 95 -17 129
rect 17 95 33 129
rect -33 79 33 95
rect -15 48 15 79
rect -15 -146 15 -120
<< polycont >>
rect -17 95 17 129
<< locali >>
rect -33 95 -17 129
rect 17 95 33 129
rect -61 36 -27 52
rect -61 -124 -27 -108
rect 27 36 61 52
rect 27 -124 61 -108
<< viali >>
rect -17 95 17 129
rect -61 -108 -27 36
rect 27 -108 61 36
<< metal1 >>
rect -29 129 29 135
rect -29 95 -17 129
rect 17 95 29 129
rect -29 89 29 95
rect -67 36 -21 48
rect -67 -108 -61 36
rect -27 -108 -21 36
rect -67 -120 -21 -108
rect 21 36 67 48
rect 21 -108 27 36
rect 61 -108 67 36
rect 21 -120 67 -108
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.84 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
