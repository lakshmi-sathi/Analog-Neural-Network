magic
tech sky130A
magscale 1 2
timestamp 1627922418
<< xpolycontact >>
rect -35 262 35 694
rect -35 -694 35 -262
<< ppolyres >>
rect -35 -262 35 262
<< viali >>
rect -19 279 19 676
rect -19 -676 19 -279
<< metal1 >>
rect -25 676 25 688
rect -25 279 -19 676
rect 19 279 25 676
rect -25 267 25 279
rect -25 -279 25 -267
rect -25 -676 -19 -279
rect 19 -676 25 -279
rect -25 -688 25 -676
<< res0p35 >>
rect -37 -264 37 264
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string parameters w 0.350 l 2.62 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 2.503k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 0.350 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
