magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_p >>
rect -1901 372 -1843 378
rect -1709 372 -1651 378
rect -1517 372 -1459 378
rect -1325 372 -1267 378
rect -1133 372 -1075 378
rect -941 372 -883 378
rect -749 372 -691 378
rect -557 372 -499 378
rect -365 372 -307 378
rect -173 372 -115 378
rect 19 372 77 378
rect 211 372 269 378
rect 403 372 461 378
rect 595 372 653 378
rect 787 372 845 378
rect 979 372 1037 378
rect 1171 372 1229 378
rect 1363 372 1421 378
rect 1555 372 1613 378
rect 1747 372 1805 378
rect 1939 372 1997 378
rect -1901 338 -1889 372
rect -1709 338 -1697 372
rect -1517 338 -1505 372
rect -1325 338 -1313 372
rect -1133 338 -1121 372
rect -941 338 -929 372
rect -749 338 -737 372
rect -557 338 -545 372
rect -365 338 -353 372
rect -173 338 -161 372
rect 19 338 31 372
rect 211 338 223 372
rect 403 338 415 372
rect 595 338 607 372
rect 787 338 799 372
rect 979 338 991 372
rect 1171 338 1183 372
rect 1363 338 1375 372
rect 1555 338 1567 372
rect 1747 338 1759 372
rect 1939 338 1951 372
rect -1901 332 -1843 338
rect -1709 332 -1651 338
rect -1517 332 -1459 338
rect -1325 332 -1267 338
rect -1133 332 -1075 338
rect -941 332 -883 338
rect -749 332 -691 338
rect -557 332 -499 338
rect -365 332 -307 338
rect -173 332 -115 338
rect 19 332 77 338
rect 211 332 269 338
rect 403 332 461 338
rect 595 332 653 338
rect 787 332 845 338
rect 979 332 1037 338
rect 1171 332 1229 338
rect 1363 332 1421 338
rect 1555 332 1613 338
rect 1747 332 1805 338
rect 1939 332 1997 338
rect -1997 -338 -1939 -332
rect -1805 -338 -1747 -332
rect -1613 -338 -1555 -332
rect -1421 -338 -1363 -332
rect -1229 -338 -1171 -332
rect -1037 -338 -979 -332
rect -845 -338 -787 -332
rect -653 -338 -595 -332
rect -461 -338 -403 -332
rect -269 -338 -211 -332
rect -77 -338 -19 -332
rect 115 -338 173 -332
rect 307 -338 365 -332
rect 499 -338 557 -332
rect 691 -338 749 -332
rect 883 -338 941 -332
rect 1075 -338 1133 -332
rect 1267 -338 1325 -332
rect 1459 -338 1517 -332
rect 1651 -338 1709 -332
rect 1843 -338 1901 -332
rect -1997 -372 -1985 -338
rect -1805 -372 -1793 -338
rect -1613 -372 -1601 -338
rect -1421 -372 -1409 -338
rect -1229 -372 -1217 -338
rect -1037 -372 -1025 -338
rect -845 -372 -833 -338
rect -653 -372 -641 -338
rect -461 -372 -449 -338
rect -269 -372 -257 -338
rect -77 -372 -65 -338
rect 115 -372 127 -338
rect 307 -372 319 -338
rect 499 -372 511 -338
rect 691 -372 703 -338
rect 883 -372 895 -338
rect 1075 -372 1087 -338
rect 1267 -372 1279 -338
rect 1459 -372 1471 -338
rect 1651 -372 1663 -338
rect 1843 -372 1855 -338
rect -1997 -378 -1939 -372
rect -1805 -378 -1747 -372
rect -1613 -378 -1555 -372
rect -1421 -378 -1363 -372
rect -1229 -378 -1171 -372
rect -1037 -378 -979 -372
rect -845 -378 -787 -372
rect -653 -378 -595 -372
rect -461 -378 -403 -372
rect -269 -378 -211 -372
rect -77 -378 -19 -372
rect 115 -378 173 -372
rect 307 -378 365 -372
rect 499 -378 557 -372
rect 691 -378 749 -372
rect 883 -378 941 -372
rect 1075 -378 1133 -372
rect 1267 -378 1325 -372
rect 1459 -378 1517 -372
rect 1651 -378 1709 -372
rect 1843 -378 1901 -372
<< pwell >>
rect -2147 440 2147 474
rect -2147 -440 -2113 440
rect 2113 -440 2147 440
rect -2147 -474 2147 -440
<< nmos >>
rect -1983 -300 -1953 300
rect -1887 -300 -1857 300
rect -1791 -300 -1761 300
rect -1695 -300 -1665 300
rect -1599 -300 -1569 300
rect -1503 -300 -1473 300
rect -1407 -300 -1377 300
rect -1311 -300 -1281 300
rect -1215 -300 -1185 300
rect -1119 -300 -1089 300
rect -1023 -300 -993 300
rect -927 -300 -897 300
rect -831 -300 -801 300
rect -735 -300 -705 300
rect -639 -300 -609 300
rect -543 -300 -513 300
rect -447 -300 -417 300
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
rect 417 -300 447 300
rect 513 -300 543 300
rect 609 -300 639 300
rect 705 -300 735 300
rect 801 -300 831 300
rect 897 -300 927 300
rect 993 -300 1023 300
rect 1089 -300 1119 300
rect 1185 -300 1215 300
rect 1281 -300 1311 300
rect 1377 -300 1407 300
rect 1473 -300 1503 300
rect 1569 -300 1599 300
rect 1665 -300 1695 300
rect 1761 -300 1791 300
rect 1857 -300 1887 300
rect 1953 -300 1983 300
<< ndiff >>
rect -2045 255 -1983 300
rect -2045 221 -2033 255
rect -1999 221 -1983 255
rect -2045 187 -1983 221
rect -2045 153 -2033 187
rect -1999 153 -1983 187
rect -2045 119 -1983 153
rect -2045 85 -2033 119
rect -1999 85 -1983 119
rect -2045 51 -1983 85
rect -2045 17 -2033 51
rect -1999 17 -1983 51
rect -2045 -17 -1983 17
rect -2045 -51 -2033 -17
rect -1999 -51 -1983 -17
rect -2045 -85 -1983 -51
rect -2045 -119 -2033 -85
rect -1999 -119 -1983 -85
rect -2045 -153 -1983 -119
rect -2045 -187 -2033 -153
rect -1999 -187 -1983 -153
rect -2045 -221 -1983 -187
rect -2045 -255 -2033 -221
rect -1999 -255 -1983 -221
rect -2045 -300 -1983 -255
rect -1953 255 -1887 300
rect -1953 221 -1937 255
rect -1903 221 -1887 255
rect -1953 187 -1887 221
rect -1953 153 -1937 187
rect -1903 153 -1887 187
rect -1953 119 -1887 153
rect -1953 85 -1937 119
rect -1903 85 -1887 119
rect -1953 51 -1887 85
rect -1953 17 -1937 51
rect -1903 17 -1887 51
rect -1953 -17 -1887 17
rect -1953 -51 -1937 -17
rect -1903 -51 -1887 -17
rect -1953 -85 -1887 -51
rect -1953 -119 -1937 -85
rect -1903 -119 -1887 -85
rect -1953 -153 -1887 -119
rect -1953 -187 -1937 -153
rect -1903 -187 -1887 -153
rect -1953 -221 -1887 -187
rect -1953 -255 -1937 -221
rect -1903 -255 -1887 -221
rect -1953 -300 -1887 -255
rect -1857 255 -1791 300
rect -1857 221 -1841 255
rect -1807 221 -1791 255
rect -1857 187 -1791 221
rect -1857 153 -1841 187
rect -1807 153 -1791 187
rect -1857 119 -1791 153
rect -1857 85 -1841 119
rect -1807 85 -1791 119
rect -1857 51 -1791 85
rect -1857 17 -1841 51
rect -1807 17 -1791 51
rect -1857 -17 -1791 17
rect -1857 -51 -1841 -17
rect -1807 -51 -1791 -17
rect -1857 -85 -1791 -51
rect -1857 -119 -1841 -85
rect -1807 -119 -1791 -85
rect -1857 -153 -1791 -119
rect -1857 -187 -1841 -153
rect -1807 -187 -1791 -153
rect -1857 -221 -1791 -187
rect -1857 -255 -1841 -221
rect -1807 -255 -1791 -221
rect -1857 -300 -1791 -255
rect -1761 255 -1695 300
rect -1761 221 -1745 255
rect -1711 221 -1695 255
rect -1761 187 -1695 221
rect -1761 153 -1745 187
rect -1711 153 -1695 187
rect -1761 119 -1695 153
rect -1761 85 -1745 119
rect -1711 85 -1695 119
rect -1761 51 -1695 85
rect -1761 17 -1745 51
rect -1711 17 -1695 51
rect -1761 -17 -1695 17
rect -1761 -51 -1745 -17
rect -1711 -51 -1695 -17
rect -1761 -85 -1695 -51
rect -1761 -119 -1745 -85
rect -1711 -119 -1695 -85
rect -1761 -153 -1695 -119
rect -1761 -187 -1745 -153
rect -1711 -187 -1695 -153
rect -1761 -221 -1695 -187
rect -1761 -255 -1745 -221
rect -1711 -255 -1695 -221
rect -1761 -300 -1695 -255
rect -1665 255 -1599 300
rect -1665 221 -1649 255
rect -1615 221 -1599 255
rect -1665 187 -1599 221
rect -1665 153 -1649 187
rect -1615 153 -1599 187
rect -1665 119 -1599 153
rect -1665 85 -1649 119
rect -1615 85 -1599 119
rect -1665 51 -1599 85
rect -1665 17 -1649 51
rect -1615 17 -1599 51
rect -1665 -17 -1599 17
rect -1665 -51 -1649 -17
rect -1615 -51 -1599 -17
rect -1665 -85 -1599 -51
rect -1665 -119 -1649 -85
rect -1615 -119 -1599 -85
rect -1665 -153 -1599 -119
rect -1665 -187 -1649 -153
rect -1615 -187 -1599 -153
rect -1665 -221 -1599 -187
rect -1665 -255 -1649 -221
rect -1615 -255 -1599 -221
rect -1665 -300 -1599 -255
rect -1569 255 -1503 300
rect -1569 221 -1553 255
rect -1519 221 -1503 255
rect -1569 187 -1503 221
rect -1569 153 -1553 187
rect -1519 153 -1503 187
rect -1569 119 -1503 153
rect -1569 85 -1553 119
rect -1519 85 -1503 119
rect -1569 51 -1503 85
rect -1569 17 -1553 51
rect -1519 17 -1503 51
rect -1569 -17 -1503 17
rect -1569 -51 -1553 -17
rect -1519 -51 -1503 -17
rect -1569 -85 -1503 -51
rect -1569 -119 -1553 -85
rect -1519 -119 -1503 -85
rect -1569 -153 -1503 -119
rect -1569 -187 -1553 -153
rect -1519 -187 -1503 -153
rect -1569 -221 -1503 -187
rect -1569 -255 -1553 -221
rect -1519 -255 -1503 -221
rect -1569 -300 -1503 -255
rect -1473 255 -1407 300
rect -1473 221 -1457 255
rect -1423 221 -1407 255
rect -1473 187 -1407 221
rect -1473 153 -1457 187
rect -1423 153 -1407 187
rect -1473 119 -1407 153
rect -1473 85 -1457 119
rect -1423 85 -1407 119
rect -1473 51 -1407 85
rect -1473 17 -1457 51
rect -1423 17 -1407 51
rect -1473 -17 -1407 17
rect -1473 -51 -1457 -17
rect -1423 -51 -1407 -17
rect -1473 -85 -1407 -51
rect -1473 -119 -1457 -85
rect -1423 -119 -1407 -85
rect -1473 -153 -1407 -119
rect -1473 -187 -1457 -153
rect -1423 -187 -1407 -153
rect -1473 -221 -1407 -187
rect -1473 -255 -1457 -221
rect -1423 -255 -1407 -221
rect -1473 -300 -1407 -255
rect -1377 255 -1311 300
rect -1377 221 -1361 255
rect -1327 221 -1311 255
rect -1377 187 -1311 221
rect -1377 153 -1361 187
rect -1327 153 -1311 187
rect -1377 119 -1311 153
rect -1377 85 -1361 119
rect -1327 85 -1311 119
rect -1377 51 -1311 85
rect -1377 17 -1361 51
rect -1327 17 -1311 51
rect -1377 -17 -1311 17
rect -1377 -51 -1361 -17
rect -1327 -51 -1311 -17
rect -1377 -85 -1311 -51
rect -1377 -119 -1361 -85
rect -1327 -119 -1311 -85
rect -1377 -153 -1311 -119
rect -1377 -187 -1361 -153
rect -1327 -187 -1311 -153
rect -1377 -221 -1311 -187
rect -1377 -255 -1361 -221
rect -1327 -255 -1311 -221
rect -1377 -300 -1311 -255
rect -1281 255 -1215 300
rect -1281 221 -1265 255
rect -1231 221 -1215 255
rect -1281 187 -1215 221
rect -1281 153 -1265 187
rect -1231 153 -1215 187
rect -1281 119 -1215 153
rect -1281 85 -1265 119
rect -1231 85 -1215 119
rect -1281 51 -1215 85
rect -1281 17 -1265 51
rect -1231 17 -1215 51
rect -1281 -17 -1215 17
rect -1281 -51 -1265 -17
rect -1231 -51 -1215 -17
rect -1281 -85 -1215 -51
rect -1281 -119 -1265 -85
rect -1231 -119 -1215 -85
rect -1281 -153 -1215 -119
rect -1281 -187 -1265 -153
rect -1231 -187 -1215 -153
rect -1281 -221 -1215 -187
rect -1281 -255 -1265 -221
rect -1231 -255 -1215 -221
rect -1281 -300 -1215 -255
rect -1185 255 -1119 300
rect -1185 221 -1169 255
rect -1135 221 -1119 255
rect -1185 187 -1119 221
rect -1185 153 -1169 187
rect -1135 153 -1119 187
rect -1185 119 -1119 153
rect -1185 85 -1169 119
rect -1135 85 -1119 119
rect -1185 51 -1119 85
rect -1185 17 -1169 51
rect -1135 17 -1119 51
rect -1185 -17 -1119 17
rect -1185 -51 -1169 -17
rect -1135 -51 -1119 -17
rect -1185 -85 -1119 -51
rect -1185 -119 -1169 -85
rect -1135 -119 -1119 -85
rect -1185 -153 -1119 -119
rect -1185 -187 -1169 -153
rect -1135 -187 -1119 -153
rect -1185 -221 -1119 -187
rect -1185 -255 -1169 -221
rect -1135 -255 -1119 -221
rect -1185 -300 -1119 -255
rect -1089 255 -1023 300
rect -1089 221 -1073 255
rect -1039 221 -1023 255
rect -1089 187 -1023 221
rect -1089 153 -1073 187
rect -1039 153 -1023 187
rect -1089 119 -1023 153
rect -1089 85 -1073 119
rect -1039 85 -1023 119
rect -1089 51 -1023 85
rect -1089 17 -1073 51
rect -1039 17 -1023 51
rect -1089 -17 -1023 17
rect -1089 -51 -1073 -17
rect -1039 -51 -1023 -17
rect -1089 -85 -1023 -51
rect -1089 -119 -1073 -85
rect -1039 -119 -1023 -85
rect -1089 -153 -1023 -119
rect -1089 -187 -1073 -153
rect -1039 -187 -1023 -153
rect -1089 -221 -1023 -187
rect -1089 -255 -1073 -221
rect -1039 -255 -1023 -221
rect -1089 -300 -1023 -255
rect -993 255 -927 300
rect -993 221 -977 255
rect -943 221 -927 255
rect -993 187 -927 221
rect -993 153 -977 187
rect -943 153 -927 187
rect -993 119 -927 153
rect -993 85 -977 119
rect -943 85 -927 119
rect -993 51 -927 85
rect -993 17 -977 51
rect -943 17 -927 51
rect -993 -17 -927 17
rect -993 -51 -977 -17
rect -943 -51 -927 -17
rect -993 -85 -927 -51
rect -993 -119 -977 -85
rect -943 -119 -927 -85
rect -993 -153 -927 -119
rect -993 -187 -977 -153
rect -943 -187 -927 -153
rect -993 -221 -927 -187
rect -993 -255 -977 -221
rect -943 -255 -927 -221
rect -993 -300 -927 -255
rect -897 255 -831 300
rect -897 221 -881 255
rect -847 221 -831 255
rect -897 187 -831 221
rect -897 153 -881 187
rect -847 153 -831 187
rect -897 119 -831 153
rect -897 85 -881 119
rect -847 85 -831 119
rect -897 51 -831 85
rect -897 17 -881 51
rect -847 17 -831 51
rect -897 -17 -831 17
rect -897 -51 -881 -17
rect -847 -51 -831 -17
rect -897 -85 -831 -51
rect -897 -119 -881 -85
rect -847 -119 -831 -85
rect -897 -153 -831 -119
rect -897 -187 -881 -153
rect -847 -187 -831 -153
rect -897 -221 -831 -187
rect -897 -255 -881 -221
rect -847 -255 -831 -221
rect -897 -300 -831 -255
rect -801 255 -735 300
rect -801 221 -785 255
rect -751 221 -735 255
rect -801 187 -735 221
rect -801 153 -785 187
rect -751 153 -735 187
rect -801 119 -735 153
rect -801 85 -785 119
rect -751 85 -735 119
rect -801 51 -735 85
rect -801 17 -785 51
rect -751 17 -735 51
rect -801 -17 -735 17
rect -801 -51 -785 -17
rect -751 -51 -735 -17
rect -801 -85 -735 -51
rect -801 -119 -785 -85
rect -751 -119 -735 -85
rect -801 -153 -735 -119
rect -801 -187 -785 -153
rect -751 -187 -735 -153
rect -801 -221 -735 -187
rect -801 -255 -785 -221
rect -751 -255 -735 -221
rect -801 -300 -735 -255
rect -705 255 -639 300
rect -705 221 -689 255
rect -655 221 -639 255
rect -705 187 -639 221
rect -705 153 -689 187
rect -655 153 -639 187
rect -705 119 -639 153
rect -705 85 -689 119
rect -655 85 -639 119
rect -705 51 -639 85
rect -705 17 -689 51
rect -655 17 -639 51
rect -705 -17 -639 17
rect -705 -51 -689 -17
rect -655 -51 -639 -17
rect -705 -85 -639 -51
rect -705 -119 -689 -85
rect -655 -119 -639 -85
rect -705 -153 -639 -119
rect -705 -187 -689 -153
rect -655 -187 -639 -153
rect -705 -221 -639 -187
rect -705 -255 -689 -221
rect -655 -255 -639 -221
rect -705 -300 -639 -255
rect -609 255 -543 300
rect -609 221 -593 255
rect -559 221 -543 255
rect -609 187 -543 221
rect -609 153 -593 187
rect -559 153 -543 187
rect -609 119 -543 153
rect -609 85 -593 119
rect -559 85 -543 119
rect -609 51 -543 85
rect -609 17 -593 51
rect -559 17 -543 51
rect -609 -17 -543 17
rect -609 -51 -593 -17
rect -559 -51 -543 -17
rect -609 -85 -543 -51
rect -609 -119 -593 -85
rect -559 -119 -543 -85
rect -609 -153 -543 -119
rect -609 -187 -593 -153
rect -559 -187 -543 -153
rect -609 -221 -543 -187
rect -609 -255 -593 -221
rect -559 -255 -543 -221
rect -609 -300 -543 -255
rect -513 255 -447 300
rect -513 221 -497 255
rect -463 221 -447 255
rect -513 187 -447 221
rect -513 153 -497 187
rect -463 153 -447 187
rect -513 119 -447 153
rect -513 85 -497 119
rect -463 85 -447 119
rect -513 51 -447 85
rect -513 17 -497 51
rect -463 17 -447 51
rect -513 -17 -447 17
rect -513 -51 -497 -17
rect -463 -51 -447 -17
rect -513 -85 -447 -51
rect -513 -119 -497 -85
rect -463 -119 -447 -85
rect -513 -153 -447 -119
rect -513 -187 -497 -153
rect -463 -187 -447 -153
rect -513 -221 -447 -187
rect -513 -255 -497 -221
rect -463 -255 -447 -221
rect -513 -300 -447 -255
rect -417 255 -351 300
rect -417 221 -401 255
rect -367 221 -351 255
rect -417 187 -351 221
rect -417 153 -401 187
rect -367 153 -351 187
rect -417 119 -351 153
rect -417 85 -401 119
rect -367 85 -351 119
rect -417 51 -351 85
rect -417 17 -401 51
rect -367 17 -351 51
rect -417 -17 -351 17
rect -417 -51 -401 -17
rect -367 -51 -351 -17
rect -417 -85 -351 -51
rect -417 -119 -401 -85
rect -367 -119 -351 -85
rect -417 -153 -351 -119
rect -417 -187 -401 -153
rect -367 -187 -351 -153
rect -417 -221 -351 -187
rect -417 -255 -401 -221
rect -367 -255 -351 -221
rect -417 -300 -351 -255
rect -321 255 -255 300
rect -321 221 -305 255
rect -271 221 -255 255
rect -321 187 -255 221
rect -321 153 -305 187
rect -271 153 -255 187
rect -321 119 -255 153
rect -321 85 -305 119
rect -271 85 -255 119
rect -321 51 -255 85
rect -321 17 -305 51
rect -271 17 -255 51
rect -321 -17 -255 17
rect -321 -51 -305 -17
rect -271 -51 -255 -17
rect -321 -85 -255 -51
rect -321 -119 -305 -85
rect -271 -119 -255 -85
rect -321 -153 -255 -119
rect -321 -187 -305 -153
rect -271 -187 -255 -153
rect -321 -221 -255 -187
rect -321 -255 -305 -221
rect -271 -255 -255 -221
rect -321 -300 -255 -255
rect -225 255 -159 300
rect -225 221 -209 255
rect -175 221 -159 255
rect -225 187 -159 221
rect -225 153 -209 187
rect -175 153 -159 187
rect -225 119 -159 153
rect -225 85 -209 119
rect -175 85 -159 119
rect -225 51 -159 85
rect -225 17 -209 51
rect -175 17 -159 51
rect -225 -17 -159 17
rect -225 -51 -209 -17
rect -175 -51 -159 -17
rect -225 -85 -159 -51
rect -225 -119 -209 -85
rect -175 -119 -159 -85
rect -225 -153 -159 -119
rect -225 -187 -209 -153
rect -175 -187 -159 -153
rect -225 -221 -159 -187
rect -225 -255 -209 -221
rect -175 -255 -159 -221
rect -225 -300 -159 -255
rect -129 255 -63 300
rect -129 221 -113 255
rect -79 221 -63 255
rect -129 187 -63 221
rect -129 153 -113 187
rect -79 153 -63 187
rect -129 119 -63 153
rect -129 85 -113 119
rect -79 85 -63 119
rect -129 51 -63 85
rect -129 17 -113 51
rect -79 17 -63 51
rect -129 -17 -63 17
rect -129 -51 -113 -17
rect -79 -51 -63 -17
rect -129 -85 -63 -51
rect -129 -119 -113 -85
rect -79 -119 -63 -85
rect -129 -153 -63 -119
rect -129 -187 -113 -153
rect -79 -187 -63 -153
rect -129 -221 -63 -187
rect -129 -255 -113 -221
rect -79 -255 -63 -221
rect -129 -300 -63 -255
rect -33 255 33 300
rect -33 221 -17 255
rect 17 221 33 255
rect -33 187 33 221
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -221 33 -187
rect -33 -255 -17 -221
rect 17 -255 33 -221
rect -33 -300 33 -255
rect 63 255 129 300
rect 63 221 79 255
rect 113 221 129 255
rect 63 187 129 221
rect 63 153 79 187
rect 113 153 129 187
rect 63 119 129 153
rect 63 85 79 119
rect 113 85 129 119
rect 63 51 129 85
rect 63 17 79 51
rect 113 17 129 51
rect 63 -17 129 17
rect 63 -51 79 -17
rect 113 -51 129 -17
rect 63 -85 129 -51
rect 63 -119 79 -85
rect 113 -119 129 -85
rect 63 -153 129 -119
rect 63 -187 79 -153
rect 113 -187 129 -153
rect 63 -221 129 -187
rect 63 -255 79 -221
rect 113 -255 129 -221
rect 63 -300 129 -255
rect 159 255 225 300
rect 159 221 175 255
rect 209 221 225 255
rect 159 187 225 221
rect 159 153 175 187
rect 209 153 225 187
rect 159 119 225 153
rect 159 85 175 119
rect 209 85 225 119
rect 159 51 225 85
rect 159 17 175 51
rect 209 17 225 51
rect 159 -17 225 17
rect 159 -51 175 -17
rect 209 -51 225 -17
rect 159 -85 225 -51
rect 159 -119 175 -85
rect 209 -119 225 -85
rect 159 -153 225 -119
rect 159 -187 175 -153
rect 209 -187 225 -153
rect 159 -221 225 -187
rect 159 -255 175 -221
rect 209 -255 225 -221
rect 159 -300 225 -255
rect 255 255 321 300
rect 255 221 271 255
rect 305 221 321 255
rect 255 187 321 221
rect 255 153 271 187
rect 305 153 321 187
rect 255 119 321 153
rect 255 85 271 119
rect 305 85 321 119
rect 255 51 321 85
rect 255 17 271 51
rect 305 17 321 51
rect 255 -17 321 17
rect 255 -51 271 -17
rect 305 -51 321 -17
rect 255 -85 321 -51
rect 255 -119 271 -85
rect 305 -119 321 -85
rect 255 -153 321 -119
rect 255 -187 271 -153
rect 305 -187 321 -153
rect 255 -221 321 -187
rect 255 -255 271 -221
rect 305 -255 321 -221
rect 255 -300 321 -255
rect 351 255 417 300
rect 351 221 367 255
rect 401 221 417 255
rect 351 187 417 221
rect 351 153 367 187
rect 401 153 417 187
rect 351 119 417 153
rect 351 85 367 119
rect 401 85 417 119
rect 351 51 417 85
rect 351 17 367 51
rect 401 17 417 51
rect 351 -17 417 17
rect 351 -51 367 -17
rect 401 -51 417 -17
rect 351 -85 417 -51
rect 351 -119 367 -85
rect 401 -119 417 -85
rect 351 -153 417 -119
rect 351 -187 367 -153
rect 401 -187 417 -153
rect 351 -221 417 -187
rect 351 -255 367 -221
rect 401 -255 417 -221
rect 351 -300 417 -255
rect 447 255 513 300
rect 447 221 463 255
rect 497 221 513 255
rect 447 187 513 221
rect 447 153 463 187
rect 497 153 513 187
rect 447 119 513 153
rect 447 85 463 119
rect 497 85 513 119
rect 447 51 513 85
rect 447 17 463 51
rect 497 17 513 51
rect 447 -17 513 17
rect 447 -51 463 -17
rect 497 -51 513 -17
rect 447 -85 513 -51
rect 447 -119 463 -85
rect 497 -119 513 -85
rect 447 -153 513 -119
rect 447 -187 463 -153
rect 497 -187 513 -153
rect 447 -221 513 -187
rect 447 -255 463 -221
rect 497 -255 513 -221
rect 447 -300 513 -255
rect 543 255 609 300
rect 543 221 559 255
rect 593 221 609 255
rect 543 187 609 221
rect 543 153 559 187
rect 593 153 609 187
rect 543 119 609 153
rect 543 85 559 119
rect 593 85 609 119
rect 543 51 609 85
rect 543 17 559 51
rect 593 17 609 51
rect 543 -17 609 17
rect 543 -51 559 -17
rect 593 -51 609 -17
rect 543 -85 609 -51
rect 543 -119 559 -85
rect 593 -119 609 -85
rect 543 -153 609 -119
rect 543 -187 559 -153
rect 593 -187 609 -153
rect 543 -221 609 -187
rect 543 -255 559 -221
rect 593 -255 609 -221
rect 543 -300 609 -255
rect 639 255 705 300
rect 639 221 655 255
rect 689 221 705 255
rect 639 187 705 221
rect 639 153 655 187
rect 689 153 705 187
rect 639 119 705 153
rect 639 85 655 119
rect 689 85 705 119
rect 639 51 705 85
rect 639 17 655 51
rect 689 17 705 51
rect 639 -17 705 17
rect 639 -51 655 -17
rect 689 -51 705 -17
rect 639 -85 705 -51
rect 639 -119 655 -85
rect 689 -119 705 -85
rect 639 -153 705 -119
rect 639 -187 655 -153
rect 689 -187 705 -153
rect 639 -221 705 -187
rect 639 -255 655 -221
rect 689 -255 705 -221
rect 639 -300 705 -255
rect 735 255 801 300
rect 735 221 751 255
rect 785 221 801 255
rect 735 187 801 221
rect 735 153 751 187
rect 785 153 801 187
rect 735 119 801 153
rect 735 85 751 119
rect 785 85 801 119
rect 735 51 801 85
rect 735 17 751 51
rect 785 17 801 51
rect 735 -17 801 17
rect 735 -51 751 -17
rect 785 -51 801 -17
rect 735 -85 801 -51
rect 735 -119 751 -85
rect 785 -119 801 -85
rect 735 -153 801 -119
rect 735 -187 751 -153
rect 785 -187 801 -153
rect 735 -221 801 -187
rect 735 -255 751 -221
rect 785 -255 801 -221
rect 735 -300 801 -255
rect 831 255 897 300
rect 831 221 847 255
rect 881 221 897 255
rect 831 187 897 221
rect 831 153 847 187
rect 881 153 897 187
rect 831 119 897 153
rect 831 85 847 119
rect 881 85 897 119
rect 831 51 897 85
rect 831 17 847 51
rect 881 17 897 51
rect 831 -17 897 17
rect 831 -51 847 -17
rect 881 -51 897 -17
rect 831 -85 897 -51
rect 831 -119 847 -85
rect 881 -119 897 -85
rect 831 -153 897 -119
rect 831 -187 847 -153
rect 881 -187 897 -153
rect 831 -221 897 -187
rect 831 -255 847 -221
rect 881 -255 897 -221
rect 831 -300 897 -255
rect 927 255 993 300
rect 927 221 943 255
rect 977 221 993 255
rect 927 187 993 221
rect 927 153 943 187
rect 977 153 993 187
rect 927 119 993 153
rect 927 85 943 119
rect 977 85 993 119
rect 927 51 993 85
rect 927 17 943 51
rect 977 17 993 51
rect 927 -17 993 17
rect 927 -51 943 -17
rect 977 -51 993 -17
rect 927 -85 993 -51
rect 927 -119 943 -85
rect 977 -119 993 -85
rect 927 -153 993 -119
rect 927 -187 943 -153
rect 977 -187 993 -153
rect 927 -221 993 -187
rect 927 -255 943 -221
rect 977 -255 993 -221
rect 927 -300 993 -255
rect 1023 255 1089 300
rect 1023 221 1039 255
rect 1073 221 1089 255
rect 1023 187 1089 221
rect 1023 153 1039 187
rect 1073 153 1089 187
rect 1023 119 1089 153
rect 1023 85 1039 119
rect 1073 85 1089 119
rect 1023 51 1089 85
rect 1023 17 1039 51
rect 1073 17 1089 51
rect 1023 -17 1089 17
rect 1023 -51 1039 -17
rect 1073 -51 1089 -17
rect 1023 -85 1089 -51
rect 1023 -119 1039 -85
rect 1073 -119 1089 -85
rect 1023 -153 1089 -119
rect 1023 -187 1039 -153
rect 1073 -187 1089 -153
rect 1023 -221 1089 -187
rect 1023 -255 1039 -221
rect 1073 -255 1089 -221
rect 1023 -300 1089 -255
rect 1119 255 1185 300
rect 1119 221 1135 255
rect 1169 221 1185 255
rect 1119 187 1185 221
rect 1119 153 1135 187
rect 1169 153 1185 187
rect 1119 119 1185 153
rect 1119 85 1135 119
rect 1169 85 1185 119
rect 1119 51 1185 85
rect 1119 17 1135 51
rect 1169 17 1185 51
rect 1119 -17 1185 17
rect 1119 -51 1135 -17
rect 1169 -51 1185 -17
rect 1119 -85 1185 -51
rect 1119 -119 1135 -85
rect 1169 -119 1185 -85
rect 1119 -153 1185 -119
rect 1119 -187 1135 -153
rect 1169 -187 1185 -153
rect 1119 -221 1185 -187
rect 1119 -255 1135 -221
rect 1169 -255 1185 -221
rect 1119 -300 1185 -255
rect 1215 255 1281 300
rect 1215 221 1231 255
rect 1265 221 1281 255
rect 1215 187 1281 221
rect 1215 153 1231 187
rect 1265 153 1281 187
rect 1215 119 1281 153
rect 1215 85 1231 119
rect 1265 85 1281 119
rect 1215 51 1281 85
rect 1215 17 1231 51
rect 1265 17 1281 51
rect 1215 -17 1281 17
rect 1215 -51 1231 -17
rect 1265 -51 1281 -17
rect 1215 -85 1281 -51
rect 1215 -119 1231 -85
rect 1265 -119 1281 -85
rect 1215 -153 1281 -119
rect 1215 -187 1231 -153
rect 1265 -187 1281 -153
rect 1215 -221 1281 -187
rect 1215 -255 1231 -221
rect 1265 -255 1281 -221
rect 1215 -300 1281 -255
rect 1311 255 1377 300
rect 1311 221 1327 255
rect 1361 221 1377 255
rect 1311 187 1377 221
rect 1311 153 1327 187
rect 1361 153 1377 187
rect 1311 119 1377 153
rect 1311 85 1327 119
rect 1361 85 1377 119
rect 1311 51 1377 85
rect 1311 17 1327 51
rect 1361 17 1377 51
rect 1311 -17 1377 17
rect 1311 -51 1327 -17
rect 1361 -51 1377 -17
rect 1311 -85 1377 -51
rect 1311 -119 1327 -85
rect 1361 -119 1377 -85
rect 1311 -153 1377 -119
rect 1311 -187 1327 -153
rect 1361 -187 1377 -153
rect 1311 -221 1377 -187
rect 1311 -255 1327 -221
rect 1361 -255 1377 -221
rect 1311 -300 1377 -255
rect 1407 255 1473 300
rect 1407 221 1423 255
rect 1457 221 1473 255
rect 1407 187 1473 221
rect 1407 153 1423 187
rect 1457 153 1473 187
rect 1407 119 1473 153
rect 1407 85 1423 119
rect 1457 85 1473 119
rect 1407 51 1473 85
rect 1407 17 1423 51
rect 1457 17 1473 51
rect 1407 -17 1473 17
rect 1407 -51 1423 -17
rect 1457 -51 1473 -17
rect 1407 -85 1473 -51
rect 1407 -119 1423 -85
rect 1457 -119 1473 -85
rect 1407 -153 1473 -119
rect 1407 -187 1423 -153
rect 1457 -187 1473 -153
rect 1407 -221 1473 -187
rect 1407 -255 1423 -221
rect 1457 -255 1473 -221
rect 1407 -300 1473 -255
rect 1503 255 1569 300
rect 1503 221 1519 255
rect 1553 221 1569 255
rect 1503 187 1569 221
rect 1503 153 1519 187
rect 1553 153 1569 187
rect 1503 119 1569 153
rect 1503 85 1519 119
rect 1553 85 1569 119
rect 1503 51 1569 85
rect 1503 17 1519 51
rect 1553 17 1569 51
rect 1503 -17 1569 17
rect 1503 -51 1519 -17
rect 1553 -51 1569 -17
rect 1503 -85 1569 -51
rect 1503 -119 1519 -85
rect 1553 -119 1569 -85
rect 1503 -153 1569 -119
rect 1503 -187 1519 -153
rect 1553 -187 1569 -153
rect 1503 -221 1569 -187
rect 1503 -255 1519 -221
rect 1553 -255 1569 -221
rect 1503 -300 1569 -255
rect 1599 255 1665 300
rect 1599 221 1615 255
rect 1649 221 1665 255
rect 1599 187 1665 221
rect 1599 153 1615 187
rect 1649 153 1665 187
rect 1599 119 1665 153
rect 1599 85 1615 119
rect 1649 85 1665 119
rect 1599 51 1665 85
rect 1599 17 1615 51
rect 1649 17 1665 51
rect 1599 -17 1665 17
rect 1599 -51 1615 -17
rect 1649 -51 1665 -17
rect 1599 -85 1665 -51
rect 1599 -119 1615 -85
rect 1649 -119 1665 -85
rect 1599 -153 1665 -119
rect 1599 -187 1615 -153
rect 1649 -187 1665 -153
rect 1599 -221 1665 -187
rect 1599 -255 1615 -221
rect 1649 -255 1665 -221
rect 1599 -300 1665 -255
rect 1695 255 1761 300
rect 1695 221 1711 255
rect 1745 221 1761 255
rect 1695 187 1761 221
rect 1695 153 1711 187
rect 1745 153 1761 187
rect 1695 119 1761 153
rect 1695 85 1711 119
rect 1745 85 1761 119
rect 1695 51 1761 85
rect 1695 17 1711 51
rect 1745 17 1761 51
rect 1695 -17 1761 17
rect 1695 -51 1711 -17
rect 1745 -51 1761 -17
rect 1695 -85 1761 -51
rect 1695 -119 1711 -85
rect 1745 -119 1761 -85
rect 1695 -153 1761 -119
rect 1695 -187 1711 -153
rect 1745 -187 1761 -153
rect 1695 -221 1761 -187
rect 1695 -255 1711 -221
rect 1745 -255 1761 -221
rect 1695 -300 1761 -255
rect 1791 255 1857 300
rect 1791 221 1807 255
rect 1841 221 1857 255
rect 1791 187 1857 221
rect 1791 153 1807 187
rect 1841 153 1857 187
rect 1791 119 1857 153
rect 1791 85 1807 119
rect 1841 85 1857 119
rect 1791 51 1857 85
rect 1791 17 1807 51
rect 1841 17 1857 51
rect 1791 -17 1857 17
rect 1791 -51 1807 -17
rect 1841 -51 1857 -17
rect 1791 -85 1857 -51
rect 1791 -119 1807 -85
rect 1841 -119 1857 -85
rect 1791 -153 1857 -119
rect 1791 -187 1807 -153
rect 1841 -187 1857 -153
rect 1791 -221 1857 -187
rect 1791 -255 1807 -221
rect 1841 -255 1857 -221
rect 1791 -300 1857 -255
rect 1887 255 1953 300
rect 1887 221 1903 255
rect 1937 221 1953 255
rect 1887 187 1953 221
rect 1887 153 1903 187
rect 1937 153 1953 187
rect 1887 119 1953 153
rect 1887 85 1903 119
rect 1937 85 1953 119
rect 1887 51 1953 85
rect 1887 17 1903 51
rect 1937 17 1953 51
rect 1887 -17 1953 17
rect 1887 -51 1903 -17
rect 1937 -51 1953 -17
rect 1887 -85 1953 -51
rect 1887 -119 1903 -85
rect 1937 -119 1953 -85
rect 1887 -153 1953 -119
rect 1887 -187 1903 -153
rect 1937 -187 1953 -153
rect 1887 -221 1953 -187
rect 1887 -255 1903 -221
rect 1937 -255 1953 -221
rect 1887 -300 1953 -255
rect 1983 255 2045 300
rect 1983 221 1999 255
rect 2033 221 2045 255
rect 1983 187 2045 221
rect 1983 153 1999 187
rect 2033 153 2045 187
rect 1983 119 2045 153
rect 1983 85 1999 119
rect 2033 85 2045 119
rect 1983 51 2045 85
rect 1983 17 1999 51
rect 2033 17 2045 51
rect 1983 -17 2045 17
rect 1983 -51 1999 -17
rect 2033 -51 2045 -17
rect 1983 -85 2045 -51
rect 1983 -119 1999 -85
rect 2033 -119 2045 -85
rect 1983 -153 2045 -119
rect 1983 -187 1999 -153
rect 2033 -187 2045 -153
rect 1983 -221 2045 -187
rect 1983 -255 1999 -221
rect 2033 -255 2045 -221
rect 1983 -300 2045 -255
<< ndiffc >>
rect -2033 221 -1999 255
rect -2033 153 -1999 187
rect -2033 85 -1999 119
rect -2033 17 -1999 51
rect -2033 -51 -1999 -17
rect -2033 -119 -1999 -85
rect -2033 -187 -1999 -153
rect -2033 -255 -1999 -221
rect -1937 221 -1903 255
rect -1937 153 -1903 187
rect -1937 85 -1903 119
rect -1937 17 -1903 51
rect -1937 -51 -1903 -17
rect -1937 -119 -1903 -85
rect -1937 -187 -1903 -153
rect -1937 -255 -1903 -221
rect -1841 221 -1807 255
rect -1841 153 -1807 187
rect -1841 85 -1807 119
rect -1841 17 -1807 51
rect -1841 -51 -1807 -17
rect -1841 -119 -1807 -85
rect -1841 -187 -1807 -153
rect -1841 -255 -1807 -221
rect -1745 221 -1711 255
rect -1745 153 -1711 187
rect -1745 85 -1711 119
rect -1745 17 -1711 51
rect -1745 -51 -1711 -17
rect -1745 -119 -1711 -85
rect -1745 -187 -1711 -153
rect -1745 -255 -1711 -221
rect -1649 221 -1615 255
rect -1649 153 -1615 187
rect -1649 85 -1615 119
rect -1649 17 -1615 51
rect -1649 -51 -1615 -17
rect -1649 -119 -1615 -85
rect -1649 -187 -1615 -153
rect -1649 -255 -1615 -221
rect -1553 221 -1519 255
rect -1553 153 -1519 187
rect -1553 85 -1519 119
rect -1553 17 -1519 51
rect -1553 -51 -1519 -17
rect -1553 -119 -1519 -85
rect -1553 -187 -1519 -153
rect -1553 -255 -1519 -221
rect -1457 221 -1423 255
rect -1457 153 -1423 187
rect -1457 85 -1423 119
rect -1457 17 -1423 51
rect -1457 -51 -1423 -17
rect -1457 -119 -1423 -85
rect -1457 -187 -1423 -153
rect -1457 -255 -1423 -221
rect -1361 221 -1327 255
rect -1361 153 -1327 187
rect -1361 85 -1327 119
rect -1361 17 -1327 51
rect -1361 -51 -1327 -17
rect -1361 -119 -1327 -85
rect -1361 -187 -1327 -153
rect -1361 -255 -1327 -221
rect -1265 221 -1231 255
rect -1265 153 -1231 187
rect -1265 85 -1231 119
rect -1265 17 -1231 51
rect -1265 -51 -1231 -17
rect -1265 -119 -1231 -85
rect -1265 -187 -1231 -153
rect -1265 -255 -1231 -221
rect -1169 221 -1135 255
rect -1169 153 -1135 187
rect -1169 85 -1135 119
rect -1169 17 -1135 51
rect -1169 -51 -1135 -17
rect -1169 -119 -1135 -85
rect -1169 -187 -1135 -153
rect -1169 -255 -1135 -221
rect -1073 221 -1039 255
rect -1073 153 -1039 187
rect -1073 85 -1039 119
rect -1073 17 -1039 51
rect -1073 -51 -1039 -17
rect -1073 -119 -1039 -85
rect -1073 -187 -1039 -153
rect -1073 -255 -1039 -221
rect -977 221 -943 255
rect -977 153 -943 187
rect -977 85 -943 119
rect -977 17 -943 51
rect -977 -51 -943 -17
rect -977 -119 -943 -85
rect -977 -187 -943 -153
rect -977 -255 -943 -221
rect -881 221 -847 255
rect -881 153 -847 187
rect -881 85 -847 119
rect -881 17 -847 51
rect -881 -51 -847 -17
rect -881 -119 -847 -85
rect -881 -187 -847 -153
rect -881 -255 -847 -221
rect -785 221 -751 255
rect -785 153 -751 187
rect -785 85 -751 119
rect -785 17 -751 51
rect -785 -51 -751 -17
rect -785 -119 -751 -85
rect -785 -187 -751 -153
rect -785 -255 -751 -221
rect -689 221 -655 255
rect -689 153 -655 187
rect -689 85 -655 119
rect -689 17 -655 51
rect -689 -51 -655 -17
rect -689 -119 -655 -85
rect -689 -187 -655 -153
rect -689 -255 -655 -221
rect -593 221 -559 255
rect -593 153 -559 187
rect -593 85 -559 119
rect -593 17 -559 51
rect -593 -51 -559 -17
rect -593 -119 -559 -85
rect -593 -187 -559 -153
rect -593 -255 -559 -221
rect -497 221 -463 255
rect -497 153 -463 187
rect -497 85 -463 119
rect -497 17 -463 51
rect -497 -51 -463 -17
rect -497 -119 -463 -85
rect -497 -187 -463 -153
rect -497 -255 -463 -221
rect -401 221 -367 255
rect -401 153 -367 187
rect -401 85 -367 119
rect -401 17 -367 51
rect -401 -51 -367 -17
rect -401 -119 -367 -85
rect -401 -187 -367 -153
rect -401 -255 -367 -221
rect -305 221 -271 255
rect -305 153 -271 187
rect -305 85 -271 119
rect -305 17 -271 51
rect -305 -51 -271 -17
rect -305 -119 -271 -85
rect -305 -187 -271 -153
rect -305 -255 -271 -221
rect -209 221 -175 255
rect -209 153 -175 187
rect -209 85 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -85
rect -209 -187 -175 -153
rect -209 -255 -175 -221
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 175 221 209 255
rect 175 153 209 187
rect 175 85 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -85
rect 175 -187 209 -153
rect 175 -255 209 -221
rect 271 221 305 255
rect 271 153 305 187
rect 271 85 305 119
rect 271 17 305 51
rect 271 -51 305 -17
rect 271 -119 305 -85
rect 271 -187 305 -153
rect 271 -255 305 -221
rect 367 221 401 255
rect 367 153 401 187
rect 367 85 401 119
rect 367 17 401 51
rect 367 -51 401 -17
rect 367 -119 401 -85
rect 367 -187 401 -153
rect 367 -255 401 -221
rect 463 221 497 255
rect 463 153 497 187
rect 463 85 497 119
rect 463 17 497 51
rect 463 -51 497 -17
rect 463 -119 497 -85
rect 463 -187 497 -153
rect 463 -255 497 -221
rect 559 221 593 255
rect 559 153 593 187
rect 559 85 593 119
rect 559 17 593 51
rect 559 -51 593 -17
rect 559 -119 593 -85
rect 559 -187 593 -153
rect 559 -255 593 -221
rect 655 221 689 255
rect 655 153 689 187
rect 655 85 689 119
rect 655 17 689 51
rect 655 -51 689 -17
rect 655 -119 689 -85
rect 655 -187 689 -153
rect 655 -255 689 -221
rect 751 221 785 255
rect 751 153 785 187
rect 751 85 785 119
rect 751 17 785 51
rect 751 -51 785 -17
rect 751 -119 785 -85
rect 751 -187 785 -153
rect 751 -255 785 -221
rect 847 221 881 255
rect 847 153 881 187
rect 847 85 881 119
rect 847 17 881 51
rect 847 -51 881 -17
rect 847 -119 881 -85
rect 847 -187 881 -153
rect 847 -255 881 -221
rect 943 221 977 255
rect 943 153 977 187
rect 943 85 977 119
rect 943 17 977 51
rect 943 -51 977 -17
rect 943 -119 977 -85
rect 943 -187 977 -153
rect 943 -255 977 -221
rect 1039 221 1073 255
rect 1039 153 1073 187
rect 1039 85 1073 119
rect 1039 17 1073 51
rect 1039 -51 1073 -17
rect 1039 -119 1073 -85
rect 1039 -187 1073 -153
rect 1039 -255 1073 -221
rect 1135 221 1169 255
rect 1135 153 1169 187
rect 1135 85 1169 119
rect 1135 17 1169 51
rect 1135 -51 1169 -17
rect 1135 -119 1169 -85
rect 1135 -187 1169 -153
rect 1135 -255 1169 -221
rect 1231 221 1265 255
rect 1231 153 1265 187
rect 1231 85 1265 119
rect 1231 17 1265 51
rect 1231 -51 1265 -17
rect 1231 -119 1265 -85
rect 1231 -187 1265 -153
rect 1231 -255 1265 -221
rect 1327 221 1361 255
rect 1327 153 1361 187
rect 1327 85 1361 119
rect 1327 17 1361 51
rect 1327 -51 1361 -17
rect 1327 -119 1361 -85
rect 1327 -187 1361 -153
rect 1327 -255 1361 -221
rect 1423 221 1457 255
rect 1423 153 1457 187
rect 1423 85 1457 119
rect 1423 17 1457 51
rect 1423 -51 1457 -17
rect 1423 -119 1457 -85
rect 1423 -187 1457 -153
rect 1423 -255 1457 -221
rect 1519 221 1553 255
rect 1519 153 1553 187
rect 1519 85 1553 119
rect 1519 17 1553 51
rect 1519 -51 1553 -17
rect 1519 -119 1553 -85
rect 1519 -187 1553 -153
rect 1519 -255 1553 -221
rect 1615 221 1649 255
rect 1615 153 1649 187
rect 1615 85 1649 119
rect 1615 17 1649 51
rect 1615 -51 1649 -17
rect 1615 -119 1649 -85
rect 1615 -187 1649 -153
rect 1615 -255 1649 -221
rect 1711 221 1745 255
rect 1711 153 1745 187
rect 1711 85 1745 119
rect 1711 17 1745 51
rect 1711 -51 1745 -17
rect 1711 -119 1745 -85
rect 1711 -187 1745 -153
rect 1711 -255 1745 -221
rect 1807 221 1841 255
rect 1807 153 1841 187
rect 1807 85 1841 119
rect 1807 17 1841 51
rect 1807 -51 1841 -17
rect 1807 -119 1841 -85
rect 1807 -187 1841 -153
rect 1807 -255 1841 -221
rect 1903 221 1937 255
rect 1903 153 1937 187
rect 1903 85 1937 119
rect 1903 17 1937 51
rect 1903 -51 1937 -17
rect 1903 -119 1937 -85
rect 1903 -187 1937 -153
rect 1903 -255 1937 -221
rect 1999 221 2033 255
rect 1999 153 2033 187
rect 1999 85 2033 119
rect 1999 17 2033 51
rect 1999 -51 2033 -17
rect 1999 -119 2033 -85
rect 1999 -187 2033 -153
rect 1999 -255 2033 -221
<< psubdiff >>
rect -2147 440 2147 474
rect -2147 357 -2113 440
rect -2147 289 -2113 323
rect 2113 357 2147 440
rect -2147 221 -2113 255
rect -2147 153 -2113 187
rect -2147 85 -2113 119
rect -2147 17 -2113 51
rect -2147 -51 -2113 -17
rect -2147 -119 -2113 -85
rect -2147 -187 -2113 -153
rect -2147 -255 -2113 -221
rect -2147 -323 -2113 -289
rect 2113 289 2147 323
rect 2113 221 2147 255
rect 2113 153 2147 187
rect 2113 85 2147 119
rect 2113 17 2147 51
rect 2113 -51 2147 -17
rect 2113 -119 2147 -85
rect 2113 -187 2147 -153
rect 2113 -255 2147 -221
rect -2147 -440 -2113 -357
rect 2113 -323 2147 -289
rect 2113 -440 2147 -357
rect -2147 -474 2147 -440
<< psubdiffcont >>
rect -2147 323 -2113 357
rect 2113 323 2147 357
rect -2147 255 -2113 289
rect -2147 187 -2113 221
rect -2147 119 -2113 153
rect -2147 51 -2113 85
rect -2147 -17 -2113 17
rect -2147 -85 -2113 -51
rect -2147 -153 -2113 -119
rect -2147 -221 -2113 -187
rect -2147 -289 -2113 -255
rect 2113 255 2147 289
rect 2113 187 2147 221
rect 2113 119 2147 153
rect 2113 51 2147 85
rect 2113 -17 2147 17
rect 2113 -85 2147 -51
rect 2113 -153 2147 -119
rect 2113 -221 2147 -187
rect 2113 -289 2147 -255
rect -2147 -357 -2113 -323
rect 2113 -357 2147 -323
<< poly >>
rect -1905 372 -1839 388
rect -1905 338 -1889 372
rect -1855 338 -1839 372
rect -1983 300 -1953 326
rect -1905 322 -1839 338
rect -1713 372 -1647 388
rect -1713 338 -1697 372
rect -1663 338 -1647 372
rect -1887 300 -1857 322
rect -1791 300 -1761 326
rect -1713 322 -1647 338
rect -1521 372 -1455 388
rect -1521 338 -1505 372
rect -1471 338 -1455 372
rect -1695 300 -1665 322
rect -1599 300 -1569 326
rect -1521 322 -1455 338
rect -1329 372 -1263 388
rect -1329 338 -1313 372
rect -1279 338 -1263 372
rect -1503 300 -1473 322
rect -1407 300 -1377 326
rect -1329 322 -1263 338
rect -1137 372 -1071 388
rect -1137 338 -1121 372
rect -1087 338 -1071 372
rect -1311 300 -1281 322
rect -1215 300 -1185 326
rect -1137 322 -1071 338
rect -945 372 -879 388
rect -945 338 -929 372
rect -895 338 -879 372
rect -1119 300 -1089 322
rect -1023 300 -993 326
rect -945 322 -879 338
rect -753 372 -687 388
rect -753 338 -737 372
rect -703 338 -687 372
rect -927 300 -897 322
rect -831 300 -801 326
rect -753 322 -687 338
rect -561 372 -495 388
rect -561 338 -545 372
rect -511 338 -495 372
rect -735 300 -705 322
rect -639 300 -609 326
rect -561 322 -495 338
rect -369 372 -303 388
rect -369 338 -353 372
rect -319 338 -303 372
rect -543 300 -513 322
rect -447 300 -417 326
rect -369 322 -303 338
rect -177 372 -111 388
rect -177 338 -161 372
rect -127 338 -111 372
rect -351 300 -321 322
rect -255 300 -225 326
rect -177 322 -111 338
rect 15 372 81 388
rect 15 338 31 372
rect 65 338 81 372
rect -159 300 -129 322
rect -63 300 -33 326
rect 15 322 81 338
rect 207 372 273 388
rect 207 338 223 372
rect 257 338 273 372
rect 33 300 63 322
rect 129 300 159 326
rect 207 322 273 338
rect 399 372 465 388
rect 399 338 415 372
rect 449 338 465 372
rect 225 300 255 322
rect 321 300 351 326
rect 399 322 465 338
rect 591 372 657 388
rect 591 338 607 372
rect 641 338 657 372
rect 417 300 447 322
rect 513 300 543 326
rect 591 322 657 338
rect 783 372 849 388
rect 783 338 799 372
rect 833 338 849 372
rect 609 300 639 322
rect 705 300 735 326
rect 783 322 849 338
rect 975 372 1041 388
rect 975 338 991 372
rect 1025 338 1041 372
rect 801 300 831 322
rect 897 300 927 326
rect 975 322 1041 338
rect 1167 372 1233 388
rect 1167 338 1183 372
rect 1217 338 1233 372
rect 993 300 1023 322
rect 1089 300 1119 326
rect 1167 322 1233 338
rect 1359 372 1425 388
rect 1359 338 1375 372
rect 1409 338 1425 372
rect 1185 300 1215 322
rect 1281 300 1311 326
rect 1359 322 1425 338
rect 1551 372 1617 388
rect 1551 338 1567 372
rect 1601 338 1617 372
rect 1377 300 1407 322
rect 1473 300 1503 326
rect 1551 322 1617 338
rect 1743 372 1809 388
rect 1743 338 1759 372
rect 1793 338 1809 372
rect 1569 300 1599 322
rect 1665 300 1695 326
rect 1743 322 1809 338
rect 1935 372 2001 388
rect 1935 338 1951 372
rect 1985 338 2001 372
rect 1761 300 1791 322
rect 1857 300 1887 326
rect 1935 322 2001 338
rect 1953 300 1983 322
rect -1983 -322 -1953 -300
rect -2001 -338 -1935 -322
rect -1887 -326 -1857 -300
rect -1791 -322 -1761 -300
rect -2001 -372 -1985 -338
rect -1951 -372 -1935 -338
rect -2001 -388 -1935 -372
rect -1809 -338 -1743 -322
rect -1695 -326 -1665 -300
rect -1599 -322 -1569 -300
rect -1809 -372 -1793 -338
rect -1759 -372 -1743 -338
rect -1809 -388 -1743 -372
rect -1617 -338 -1551 -322
rect -1503 -326 -1473 -300
rect -1407 -322 -1377 -300
rect -1617 -372 -1601 -338
rect -1567 -372 -1551 -338
rect -1617 -388 -1551 -372
rect -1425 -338 -1359 -322
rect -1311 -326 -1281 -300
rect -1215 -322 -1185 -300
rect -1425 -372 -1409 -338
rect -1375 -372 -1359 -338
rect -1425 -388 -1359 -372
rect -1233 -338 -1167 -322
rect -1119 -326 -1089 -300
rect -1023 -322 -993 -300
rect -1233 -372 -1217 -338
rect -1183 -372 -1167 -338
rect -1233 -388 -1167 -372
rect -1041 -338 -975 -322
rect -927 -326 -897 -300
rect -831 -322 -801 -300
rect -1041 -372 -1025 -338
rect -991 -372 -975 -338
rect -1041 -388 -975 -372
rect -849 -338 -783 -322
rect -735 -326 -705 -300
rect -639 -322 -609 -300
rect -849 -372 -833 -338
rect -799 -372 -783 -338
rect -849 -388 -783 -372
rect -657 -338 -591 -322
rect -543 -326 -513 -300
rect -447 -322 -417 -300
rect -657 -372 -641 -338
rect -607 -372 -591 -338
rect -657 -388 -591 -372
rect -465 -338 -399 -322
rect -351 -326 -321 -300
rect -255 -322 -225 -300
rect -465 -372 -449 -338
rect -415 -372 -399 -338
rect -465 -388 -399 -372
rect -273 -338 -207 -322
rect -159 -326 -129 -300
rect -63 -322 -33 -300
rect -273 -372 -257 -338
rect -223 -372 -207 -338
rect -273 -388 -207 -372
rect -81 -338 -15 -322
rect 33 -326 63 -300
rect 129 -322 159 -300
rect -81 -372 -65 -338
rect -31 -372 -15 -338
rect -81 -388 -15 -372
rect 111 -338 177 -322
rect 225 -326 255 -300
rect 321 -322 351 -300
rect 111 -372 127 -338
rect 161 -372 177 -338
rect 111 -388 177 -372
rect 303 -338 369 -322
rect 417 -326 447 -300
rect 513 -322 543 -300
rect 303 -372 319 -338
rect 353 -372 369 -338
rect 303 -388 369 -372
rect 495 -338 561 -322
rect 609 -326 639 -300
rect 705 -322 735 -300
rect 495 -372 511 -338
rect 545 -372 561 -338
rect 495 -388 561 -372
rect 687 -338 753 -322
rect 801 -326 831 -300
rect 897 -322 927 -300
rect 687 -372 703 -338
rect 737 -372 753 -338
rect 687 -388 753 -372
rect 879 -338 945 -322
rect 993 -326 1023 -300
rect 1089 -322 1119 -300
rect 879 -372 895 -338
rect 929 -372 945 -338
rect 879 -388 945 -372
rect 1071 -338 1137 -322
rect 1185 -326 1215 -300
rect 1281 -322 1311 -300
rect 1071 -372 1087 -338
rect 1121 -372 1137 -338
rect 1071 -388 1137 -372
rect 1263 -338 1329 -322
rect 1377 -326 1407 -300
rect 1473 -322 1503 -300
rect 1263 -372 1279 -338
rect 1313 -372 1329 -338
rect 1263 -388 1329 -372
rect 1455 -338 1521 -322
rect 1569 -326 1599 -300
rect 1665 -322 1695 -300
rect 1455 -372 1471 -338
rect 1505 -372 1521 -338
rect 1455 -388 1521 -372
rect 1647 -338 1713 -322
rect 1761 -326 1791 -300
rect 1857 -322 1887 -300
rect 1647 -372 1663 -338
rect 1697 -372 1713 -338
rect 1647 -388 1713 -372
rect 1839 -338 1905 -322
rect 1953 -326 1983 -300
rect 1839 -372 1855 -338
rect 1889 -372 1905 -338
rect 1839 -388 1905 -372
<< polycont >>
rect -1889 338 -1855 372
rect -1697 338 -1663 372
rect -1505 338 -1471 372
rect -1313 338 -1279 372
rect -1121 338 -1087 372
rect -929 338 -895 372
rect -737 338 -703 372
rect -545 338 -511 372
rect -353 338 -319 372
rect -161 338 -127 372
rect 31 338 65 372
rect 223 338 257 372
rect 415 338 449 372
rect 607 338 641 372
rect 799 338 833 372
rect 991 338 1025 372
rect 1183 338 1217 372
rect 1375 338 1409 372
rect 1567 338 1601 372
rect 1759 338 1793 372
rect 1951 338 1985 372
rect -1985 -372 -1951 -338
rect -1793 -372 -1759 -338
rect -1601 -372 -1567 -338
rect -1409 -372 -1375 -338
rect -1217 -372 -1183 -338
rect -1025 -372 -991 -338
rect -833 -372 -799 -338
rect -641 -372 -607 -338
rect -449 -372 -415 -338
rect -257 -372 -223 -338
rect -65 -372 -31 -338
rect 127 -372 161 -338
rect 319 -372 353 -338
rect 511 -372 545 -338
rect 703 -372 737 -338
rect 895 -372 929 -338
rect 1087 -372 1121 -338
rect 1279 -372 1313 -338
rect 1471 -372 1505 -338
rect 1663 -372 1697 -338
rect 1855 -372 1889 -338
<< locali >>
rect -2147 440 2147 474
rect -2147 357 -2113 440
rect -1905 338 -1889 372
rect -1855 338 -1839 372
rect -1713 338 -1697 372
rect -1663 338 -1647 372
rect -1521 338 -1505 372
rect -1471 338 -1455 372
rect -1329 338 -1313 372
rect -1279 338 -1263 372
rect -1137 338 -1121 372
rect -1087 338 -1071 372
rect -945 338 -929 372
rect -895 338 -879 372
rect -753 338 -737 372
rect -703 338 -687 372
rect -561 338 -545 372
rect -511 338 -495 372
rect -369 338 -353 372
rect -319 338 -303 372
rect -177 338 -161 372
rect -127 338 -111 372
rect 15 338 31 372
rect 65 338 81 372
rect 207 338 223 372
rect 257 338 273 372
rect 399 338 415 372
rect 449 338 465 372
rect 591 338 607 372
rect 641 338 657 372
rect 783 338 799 372
rect 833 338 849 372
rect 975 338 991 372
rect 1025 338 1041 372
rect 1167 338 1183 372
rect 1217 338 1233 372
rect 1359 338 1375 372
rect 1409 338 1425 372
rect 1551 338 1567 372
rect 1601 338 1617 372
rect 1743 338 1759 372
rect 1793 338 1809 372
rect 1935 338 1951 372
rect 1985 338 2001 372
rect 2113 357 2147 440
rect -2147 289 -2113 323
rect -2147 221 -2113 255
rect -2147 153 -2113 187
rect -2147 85 -2113 119
rect -2147 17 -2113 51
rect -2147 -51 -2113 -17
rect -2147 -119 -2113 -85
rect -2147 -187 -2113 -153
rect -2147 -255 -2113 -221
rect -2147 -323 -2113 -289
rect -2033 269 -1999 304
rect -2033 197 -1999 221
rect -2033 125 -1999 153
rect -2033 53 -1999 85
rect -2033 -17 -1999 17
rect -2033 -85 -1999 -53
rect -2033 -153 -1999 -125
rect -2033 -221 -1999 -197
rect -2033 -304 -1999 -269
rect -1937 269 -1903 304
rect -1937 197 -1903 221
rect -1937 125 -1903 153
rect -1937 53 -1903 85
rect -1937 -17 -1903 17
rect -1937 -85 -1903 -53
rect -1937 -153 -1903 -125
rect -1937 -221 -1903 -197
rect -1937 -304 -1903 -269
rect -1841 269 -1807 304
rect -1841 197 -1807 221
rect -1841 125 -1807 153
rect -1841 53 -1807 85
rect -1841 -17 -1807 17
rect -1841 -85 -1807 -53
rect -1841 -153 -1807 -125
rect -1841 -221 -1807 -197
rect -1841 -304 -1807 -269
rect -1745 269 -1711 304
rect -1745 197 -1711 221
rect -1745 125 -1711 153
rect -1745 53 -1711 85
rect -1745 -17 -1711 17
rect -1745 -85 -1711 -53
rect -1745 -153 -1711 -125
rect -1745 -221 -1711 -197
rect -1745 -304 -1711 -269
rect -1649 269 -1615 304
rect -1649 197 -1615 221
rect -1649 125 -1615 153
rect -1649 53 -1615 85
rect -1649 -17 -1615 17
rect -1649 -85 -1615 -53
rect -1649 -153 -1615 -125
rect -1649 -221 -1615 -197
rect -1649 -304 -1615 -269
rect -1553 269 -1519 304
rect -1553 197 -1519 221
rect -1553 125 -1519 153
rect -1553 53 -1519 85
rect -1553 -17 -1519 17
rect -1553 -85 -1519 -53
rect -1553 -153 -1519 -125
rect -1553 -221 -1519 -197
rect -1553 -304 -1519 -269
rect -1457 269 -1423 304
rect -1457 197 -1423 221
rect -1457 125 -1423 153
rect -1457 53 -1423 85
rect -1457 -17 -1423 17
rect -1457 -85 -1423 -53
rect -1457 -153 -1423 -125
rect -1457 -221 -1423 -197
rect -1457 -304 -1423 -269
rect -1361 269 -1327 304
rect -1361 197 -1327 221
rect -1361 125 -1327 153
rect -1361 53 -1327 85
rect -1361 -17 -1327 17
rect -1361 -85 -1327 -53
rect -1361 -153 -1327 -125
rect -1361 -221 -1327 -197
rect -1361 -304 -1327 -269
rect -1265 269 -1231 304
rect -1265 197 -1231 221
rect -1265 125 -1231 153
rect -1265 53 -1231 85
rect -1265 -17 -1231 17
rect -1265 -85 -1231 -53
rect -1265 -153 -1231 -125
rect -1265 -221 -1231 -197
rect -1265 -304 -1231 -269
rect -1169 269 -1135 304
rect -1169 197 -1135 221
rect -1169 125 -1135 153
rect -1169 53 -1135 85
rect -1169 -17 -1135 17
rect -1169 -85 -1135 -53
rect -1169 -153 -1135 -125
rect -1169 -221 -1135 -197
rect -1169 -304 -1135 -269
rect -1073 269 -1039 304
rect -1073 197 -1039 221
rect -1073 125 -1039 153
rect -1073 53 -1039 85
rect -1073 -17 -1039 17
rect -1073 -85 -1039 -53
rect -1073 -153 -1039 -125
rect -1073 -221 -1039 -197
rect -1073 -304 -1039 -269
rect -977 269 -943 304
rect -977 197 -943 221
rect -977 125 -943 153
rect -977 53 -943 85
rect -977 -17 -943 17
rect -977 -85 -943 -53
rect -977 -153 -943 -125
rect -977 -221 -943 -197
rect -977 -304 -943 -269
rect -881 269 -847 304
rect -881 197 -847 221
rect -881 125 -847 153
rect -881 53 -847 85
rect -881 -17 -847 17
rect -881 -85 -847 -53
rect -881 -153 -847 -125
rect -881 -221 -847 -197
rect -881 -304 -847 -269
rect -785 269 -751 304
rect -785 197 -751 221
rect -785 125 -751 153
rect -785 53 -751 85
rect -785 -17 -751 17
rect -785 -85 -751 -53
rect -785 -153 -751 -125
rect -785 -221 -751 -197
rect -785 -304 -751 -269
rect -689 269 -655 304
rect -689 197 -655 221
rect -689 125 -655 153
rect -689 53 -655 85
rect -689 -17 -655 17
rect -689 -85 -655 -53
rect -689 -153 -655 -125
rect -689 -221 -655 -197
rect -689 -304 -655 -269
rect -593 269 -559 304
rect -593 197 -559 221
rect -593 125 -559 153
rect -593 53 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -53
rect -593 -153 -559 -125
rect -593 -221 -559 -197
rect -593 -304 -559 -269
rect -497 269 -463 304
rect -497 197 -463 221
rect -497 125 -463 153
rect -497 53 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -53
rect -497 -153 -463 -125
rect -497 -221 -463 -197
rect -497 -304 -463 -269
rect -401 269 -367 304
rect -401 197 -367 221
rect -401 125 -367 153
rect -401 53 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -53
rect -401 -153 -367 -125
rect -401 -221 -367 -197
rect -401 -304 -367 -269
rect -305 269 -271 304
rect -305 197 -271 221
rect -305 125 -271 153
rect -305 53 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -53
rect -305 -153 -271 -125
rect -305 -221 -271 -197
rect -305 -304 -271 -269
rect -209 269 -175 304
rect -209 197 -175 221
rect -209 125 -175 153
rect -209 53 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -53
rect -209 -153 -175 -125
rect -209 -221 -175 -197
rect -209 -304 -175 -269
rect -113 269 -79 304
rect -113 197 -79 221
rect -113 125 -79 153
rect -113 53 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -53
rect -113 -153 -79 -125
rect -113 -221 -79 -197
rect -113 -304 -79 -269
rect -17 269 17 304
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -304 17 -269
rect 79 269 113 304
rect 79 197 113 221
rect 79 125 113 153
rect 79 53 113 85
rect 79 -17 113 17
rect 79 -85 113 -53
rect 79 -153 113 -125
rect 79 -221 113 -197
rect 79 -304 113 -269
rect 175 269 209 304
rect 175 197 209 221
rect 175 125 209 153
rect 175 53 209 85
rect 175 -17 209 17
rect 175 -85 209 -53
rect 175 -153 209 -125
rect 175 -221 209 -197
rect 175 -304 209 -269
rect 271 269 305 304
rect 271 197 305 221
rect 271 125 305 153
rect 271 53 305 85
rect 271 -17 305 17
rect 271 -85 305 -53
rect 271 -153 305 -125
rect 271 -221 305 -197
rect 271 -304 305 -269
rect 367 269 401 304
rect 367 197 401 221
rect 367 125 401 153
rect 367 53 401 85
rect 367 -17 401 17
rect 367 -85 401 -53
rect 367 -153 401 -125
rect 367 -221 401 -197
rect 367 -304 401 -269
rect 463 269 497 304
rect 463 197 497 221
rect 463 125 497 153
rect 463 53 497 85
rect 463 -17 497 17
rect 463 -85 497 -53
rect 463 -153 497 -125
rect 463 -221 497 -197
rect 463 -304 497 -269
rect 559 269 593 304
rect 559 197 593 221
rect 559 125 593 153
rect 559 53 593 85
rect 559 -17 593 17
rect 559 -85 593 -53
rect 559 -153 593 -125
rect 559 -221 593 -197
rect 559 -304 593 -269
rect 655 269 689 304
rect 655 197 689 221
rect 655 125 689 153
rect 655 53 689 85
rect 655 -17 689 17
rect 655 -85 689 -53
rect 655 -153 689 -125
rect 655 -221 689 -197
rect 655 -304 689 -269
rect 751 269 785 304
rect 751 197 785 221
rect 751 125 785 153
rect 751 53 785 85
rect 751 -17 785 17
rect 751 -85 785 -53
rect 751 -153 785 -125
rect 751 -221 785 -197
rect 751 -304 785 -269
rect 847 269 881 304
rect 847 197 881 221
rect 847 125 881 153
rect 847 53 881 85
rect 847 -17 881 17
rect 847 -85 881 -53
rect 847 -153 881 -125
rect 847 -221 881 -197
rect 847 -304 881 -269
rect 943 269 977 304
rect 943 197 977 221
rect 943 125 977 153
rect 943 53 977 85
rect 943 -17 977 17
rect 943 -85 977 -53
rect 943 -153 977 -125
rect 943 -221 977 -197
rect 943 -304 977 -269
rect 1039 269 1073 304
rect 1039 197 1073 221
rect 1039 125 1073 153
rect 1039 53 1073 85
rect 1039 -17 1073 17
rect 1039 -85 1073 -53
rect 1039 -153 1073 -125
rect 1039 -221 1073 -197
rect 1039 -304 1073 -269
rect 1135 269 1169 304
rect 1135 197 1169 221
rect 1135 125 1169 153
rect 1135 53 1169 85
rect 1135 -17 1169 17
rect 1135 -85 1169 -53
rect 1135 -153 1169 -125
rect 1135 -221 1169 -197
rect 1135 -304 1169 -269
rect 1231 269 1265 304
rect 1231 197 1265 221
rect 1231 125 1265 153
rect 1231 53 1265 85
rect 1231 -17 1265 17
rect 1231 -85 1265 -53
rect 1231 -153 1265 -125
rect 1231 -221 1265 -197
rect 1231 -304 1265 -269
rect 1327 269 1361 304
rect 1327 197 1361 221
rect 1327 125 1361 153
rect 1327 53 1361 85
rect 1327 -17 1361 17
rect 1327 -85 1361 -53
rect 1327 -153 1361 -125
rect 1327 -221 1361 -197
rect 1327 -304 1361 -269
rect 1423 269 1457 304
rect 1423 197 1457 221
rect 1423 125 1457 153
rect 1423 53 1457 85
rect 1423 -17 1457 17
rect 1423 -85 1457 -53
rect 1423 -153 1457 -125
rect 1423 -221 1457 -197
rect 1423 -304 1457 -269
rect 1519 269 1553 304
rect 1519 197 1553 221
rect 1519 125 1553 153
rect 1519 53 1553 85
rect 1519 -17 1553 17
rect 1519 -85 1553 -53
rect 1519 -153 1553 -125
rect 1519 -221 1553 -197
rect 1519 -304 1553 -269
rect 1615 269 1649 304
rect 1615 197 1649 221
rect 1615 125 1649 153
rect 1615 53 1649 85
rect 1615 -17 1649 17
rect 1615 -85 1649 -53
rect 1615 -153 1649 -125
rect 1615 -221 1649 -197
rect 1615 -304 1649 -269
rect 1711 269 1745 304
rect 1711 197 1745 221
rect 1711 125 1745 153
rect 1711 53 1745 85
rect 1711 -17 1745 17
rect 1711 -85 1745 -53
rect 1711 -153 1745 -125
rect 1711 -221 1745 -197
rect 1711 -304 1745 -269
rect 1807 269 1841 304
rect 1807 197 1841 221
rect 1807 125 1841 153
rect 1807 53 1841 85
rect 1807 -17 1841 17
rect 1807 -85 1841 -53
rect 1807 -153 1841 -125
rect 1807 -221 1841 -197
rect 1807 -304 1841 -269
rect 1903 269 1937 304
rect 1903 197 1937 221
rect 1903 125 1937 153
rect 1903 53 1937 85
rect 1903 -17 1937 17
rect 1903 -85 1937 -53
rect 1903 -153 1937 -125
rect 1903 -221 1937 -197
rect 1903 -304 1937 -269
rect 1999 269 2033 304
rect 1999 197 2033 221
rect 1999 125 2033 153
rect 1999 53 2033 85
rect 1999 -17 2033 17
rect 1999 -85 2033 -53
rect 1999 -153 2033 -125
rect 1999 -221 2033 -197
rect 1999 -304 2033 -269
rect 2113 289 2147 323
rect 2113 221 2147 255
rect 2113 153 2147 187
rect 2113 85 2147 119
rect 2113 17 2147 51
rect 2113 -51 2147 -17
rect 2113 -119 2147 -85
rect 2113 -187 2147 -153
rect 2113 -255 2147 -221
rect 2113 -323 2147 -289
rect -2147 -440 -2113 -357
rect -2001 -372 -1985 -338
rect -1951 -372 -1935 -338
rect -1809 -372 -1793 -338
rect -1759 -372 -1743 -338
rect -1617 -372 -1601 -338
rect -1567 -372 -1551 -338
rect -1425 -372 -1409 -338
rect -1375 -372 -1359 -338
rect -1233 -372 -1217 -338
rect -1183 -372 -1167 -338
rect -1041 -372 -1025 -338
rect -991 -372 -975 -338
rect -849 -372 -833 -338
rect -799 -372 -783 -338
rect -657 -372 -641 -338
rect -607 -372 -591 -338
rect -465 -372 -449 -338
rect -415 -372 -399 -338
rect -273 -372 -257 -338
rect -223 -372 -207 -338
rect -81 -372 -65 -338
rect -31 -372 -15 -338
rect 111 -372 127 -338
rect 161 -372 177 -338
rect 303 -372 319 -338
rect 353 -372 369 -338
rect 495 -372 511 -338
rect 545 -372 561 -338
rect 687 -372 703 -338
rect 737 -372 753 -338
rect 879 -372 895 -338
rect 929 -372 945 -338
rect 1071 -372 1087 -338
rect 1121 -372 1137 -338
rect 1263 -372 1279 -338
rect 1313 -372 1329 -338
rect 1455 -372 1471 -338
rect 1505 -372 1521 -338
rect 1647 -372 1663 -338
rect 1697 -372 1713 -338
rect 1839 -372 1855 -338
rect 1889 -372 1905 -338
rect 2113 -440 2147 -357
rect -2147 -474 2147 -440
<< viali >>
rect -1889 338 -1855 372
rect -1697 338 -1663 372
rect -1505 338 -1471 372
rect -1313 338 -1279 372
rect -1121 338 -1087 372
rect -929 338 -895 372
rect -737 338 -703 372
rect -545 338 -511 372
rect -353 338 -319 372
rect -161 338 -127 372
rect 31 338 65 372
rect 223 338 257 372
rect 415 338 449 372
rect 607 338 641 372
rect 799 338 833 372
rect 991 338 1025 372
rect 1183 338 1217 372
rect 1375 338 1409 372
rect 1567 338 1601 372
rect 1759 338 1793 372
rect 1951 338 1985 372
rect -2033 255 -1999 269
rect -2033 235 -1999 255
rect -2033 187 -1999 197
rect -2033 163 -1999 187
rect -2033 119 -1999 125
rect -2033 91 -1999 119
rect -2033 51 -1999 53
rect -2033 19 -1999 51
rect -2033 -51 -1999 -19
rect -2033 -53 -1999 -51
rect -2033 -119 -1999 -91
rect -2033 -125 -1999 -119
rect -2033 -187 -1999 -163
rect -2033 -197 -1999 -187
rect -2033 -255 -1999 -235
rect -2033 -269 -1999 -255
rect -1937 255 -1903 269
rect -1937 235 -1903 255
rect -1937 187 -1903 197
rect -1937 163 -1903 187
rect -1937 119 -1903 125
rect -1937 91 -1903 119
rect -1937 51 -1903 53
rect -1937 19 -1903 51
rect -1937 -51 -1903 -19
rect -1937 -53 -1903 -51
rect -1937 -119 -1903 -91
rect -1937 -125 -1903 -119
rect -1937 -187 -1903 -163
rect -1937 -197 -1903 -187
rect -1937 -255 -1903 -235
rect -1937 -269 -1903 -255
rect -1841 255 -1807 269
rect -1841 235 -1807 255
rect -1841 187 -1807 197
rect -1841 163 -1807 187
rect -1841 119 -1807 125
rect -1841 91 -1807 119
rect -1841 51 -1807 53
rect -1841 19 -1807 51
rect -1841 -51 -1807 -19
rect -1841 -53 -1807 -51
rect -1841 -119 -1807 -91
rect -1841 -125 -1807 -119
rect -1841 -187 -1807 -163
rect -1841 -197 -1807 -187
rect -1841 -255 -1807 -235
rect -1841 -269 -1807 -255
rect -1745 255 -1711 269
rect -1745 235 -1711 255
rect -1745 187 -1711 197
rect -1745 163 -1711 187
rect -1745 119 -1711 125
rect -1745 91 -1711 119
rect -1745 51 -1711 53
rect -1745 19 -1711 51
rect -1745 -51 -1711 -19
rect -1745 -53 -1711 -51
rect -1745 -119 -1711 -91
rect -1745 -125 -1711 -119
rect -1745 -187 -1711 -163
rect -1745 -197 -1711 -187
rect -1745 -255 -1711 -235
rect -1745 -269 -1711 -255
rect -1649 255 -1615 269
rect -1649 235 -1615 255
rect -1649 187 -1615 197
rect -1649 163 -1615 187
rect -1649 119 -1615 125
rect -1649 91 -1615 119
rect -1649 51 -1615 53
rect -1649 19 -1615 51
rect -1649 -51 -1615 -19
rect -1649 -53 -1615 -51
rect -1649 -119 -1615 -91
rect -1649 -125 -1615 -119
rect -1649 -187 -1615 -163
rect -1649 -197 -1615 -187
rect -1649 -255 -1615 -235
rect -1649 -269 -1615 -255
rect -1553 255 -1519 269
rect -1553 235 -1519 255
rect -1553 187 -1519 197
rect -1553 163 -1519 187
rect -1553 119 -1519 125
rect -1553 91 -1519 119
rect -1553 51 -1519 53
rect -1553 19 -1519 51
rect -1553 -51 -1519 -19
rect -1553 -53 -1519 -51
rect -1553 -119 -1519 -91
rect -1553 -125 -1519 -119
rect -1553 -187 -1519 -163
rect -1553 -197 -1519 -187
rect -1553 -255 -1519 -235
rect -1553 -269 -1519 -255
rect -1457 255 -1423 269
rect -1457 235 -1423 255
rect -1457 187 -1423 197
rect -1457 163 -1423 187
rect -1457 119 -1423 125
rect -1457 91 -1423 119
rect -1457 51 -1423 53
rect -1457 19 -1423 51
rect -1457 -51 -1423 -19
rect -1457 -53 -1423 -51
rect -1457 -119 -1423 -91
rect -1457 -125 -1423 -119
rect -1457 -187 -1423 -163
rect -1457 -197 -1423 -187
rect -1457 -255 -1423 -235
rect -1457 -269 -1423 -255
rect -1361 255 -1327 269
rect -1361 235 -1327 255
rect -1361 187 -1327 197
rect -1361 163 -1327 187
rect -1361 119 -1327 125
rect -1361 91 -1327 119
rect -1361 51 -1327 53
rect -1361 19 -1327 51
rect -1361 -51 -1327 -19
rect -1361 -53 -1327 -51
rect -1361 -119 -1327 -91
rect -1361 -125 -1327 -119
rect -1361 -187 -1327 -163
rect -1361 -197 -1327 -187
rect -1361 -255 -1327 -235
rect -1361 -269 -1327 -255
rect -1265 255 -1231 269
rect -1265 235 -1231 255
rect -1265 187 -1231 197
rect -1265 163 -1231 187
rect -1265 119 -1231 125
rect -1265 91 -1231 119
rect -1265 51 -1231 53
rect -1265 19 -1231 51
rect -1265 -51 -1231 -19
rect -1265 -53 -1231 -51
rect -1265 -119 -1231 -91
rect -1265 -125 -1231 -119
rect -1265 -187 -1231 -163
rect -1265 -197 -1231 -187
rect -1265 -255 -1231 -235
rect -1265 -269 -1231 -255
rect -1169 255 -1135 269
rect -1169 235 -1135 255
rect -1169 187 -1135 197
rect -1169 163 -1135 187
rect -1169 119 -1135 125
rect -1169 91 -1135 119
rect -1169 51 -1135 53
rect -1169 19 -1135 51
rect -1169 -51 -1135 -19
rect -1169 -53 -1135 -51
rect -1169 -119 -1135 -91
rect -1169 -125 -1135 -119
rect -1169 -187 -1135 -163
rect -1169 -197 -1135 -187
rect -1169 -255 -1135 -235
rect -1169 -269 -1135 -255
rect -1073 255 -1039 269
rect -1073 235 -1039 255
rect -1073 187 -1039 197
rect -1073 163 -1039 187
rect -1073 119 -1039 125
rect -1073 91 -1039 119
rect -1073 51 -1039 53
rect -1073 19 -1039 51
rect -1073 -51 -1039 -19
rect -1073 -53 -1039 -51
rect -1073 -119 -1039 -91
rect -1073 -125 -1039 -119
rect -1073 -187 -1039 -163
rect -1073 -197 -1039 -187
rect -1073 -255 -1039 -235
rect -1073 -269 -1039 -255
rect -977 255 -943 269
rect -977 235 -943 255
rect -977 187 -943 197
rect -977 163 -943 187
rect -977 119 -943 125
rect -977 91 -943 119
rect -977 51 -943 53
rect -977 19 -943 51
rect -977 -51 -943 -19
rect -977 -53 -943 -51
rect -977 -119 -943 -91
rect -977 -125 -943 -119
rect -977 -187 -943 -163
rect -977 -197 -943 -187
rect -977 -255 -943 -235
rect -977 -269 -943 -255
rect -881 255 -847 269
rect -881 235 -847 255
rect -881 187 -847 197
rect -881 163 -847 187
rect -881 119 -847 125
rect -881 91 -847 119
rect -881 51 -847 53
rect -881 19 -847 51
rect -881 -51 -847 -19
rect -881 -53 -847 -51
rect -881 -119 -847 -91
rect -881 -125 -847 -119
rect -881 -187 -847 -163
rect -881 -197 -847 -187
rect -881 -255 -847 -235
rect -881 -269 -847 -255
rect -785 255 -751 269
rect -785 235 -751 255
rect -785 187 -751 197
rect -785 163 -751 187
rect -785 119 -751 125
rect -785 91 -751 119
rect -785 51 -751 53
rect -785 19 -751 51
rect -785 -51 -751 -19
rect -785 -53 -751 -51
rect -785 -119 -751 -91
rect -785 -125 -751 -119
rect -785 -187 -751 -163
rect -785 -197 -751 -187
rect -785 -255 -751 -235
rect -785 -269 -751 -255
rect -689 255 -655 269
rect -689 235 -655 255
rect -689 187 -655 197
rect -689 163 -655 187
rect -689 119 -655 125
rect -689 91 -655 119
rect -689 51 -655 53
rect -689 19 -655 51
rect -689 -51 -655 -19
rect -689 -53 -655 -51
rect -689 -119 -655 -91
rect -689 -125 -655 -119
rect -689 -187 -655 -163
rect -689 -197 -655 -187
rect -689 -255 -655 -235
rect -689 -269 -655 -255
rect -593 255 -559 269
rect -593 235 -559 255
rect -593 187 -559 197
rect -593 163 -559 187
rect -593 119 -559 125
rect -593 91 -559 119
rect -593 51 -559 53
rect -593 19 -559 51
rect -593 -51 -559 -19
rect -593 -53 -559 -51
rect -593 -119 -559 -91
rect -593 -125 -559 -119
rect -593 -187 -559 -163
rect -593 -197 -559 -187
rect -593 -255 -559 -235
rect -593 -269 -559 -255
rect -497 255 -463 269
rect -497 235 -463 255
rect -497 187 -463 197
rect -497 163 -463 187
rect -497 119 -463 125
rect -497 91 -463 119
rect -497 51 -463 53
rect -497 19 -463 51
rect -497 -51 -463 -19
rect -497 -53 -463 -51
rect -497 -119 -463 -91
rect -497 -125 -463 -119
rect -497 -187 -463 -163
rect -497 -197 -463 -187
rect -497 -255 -463 -235
rect -497 -269 -463 -255
rect -401 255 -367 269
rect -401 235 -367 255
rect -401 187 -367 197
rect -401 163 -367 187
rect -401 119 -367 125
rect -401 91 -367 119
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -401 -119 -367 -91
rect -401 -125 -367 -119
rect -401 -187 -367 -163
rect -401 -197 -367 -187
rect -401 -255 -367 -235
rect -401 -269 -367 -255
rect -305 255 -271 269
rect -305 235 -271 255
rect -305 187 -271 197
rect -305 163 -271 187
rect -305 119 -271 125
rect -305 91 -271 119
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -305 -119 -271 -91
rect -305 -125 -271 -119
rect -305 -187 -271 -163
rect -305 -197 -271 -187
rect -305 -255 -271 -235
rect -305 -269 -271 -255
rect -209 255 -175 269
rect -209 235 -175 255
rect -209 187 -175 197
rect -209 163 -175 187
rect -209 119 -175 125
rect -209 91 -175 119
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -209 -119 -175 -91
rect -209 -125 -175 -119
rect -209 -187 -175 -163
rect -209 -197 -175 -187
rect -209 -255 -175 -235
rect -209 -269 -175 -255
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 175 255 209 269
rect 175 235 209 255
rect 175 187 209 197
rect 175 163 209 187
rect 175 119 209 125
rect 175 91 209 119
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 175 -119 209 -91
rect 175 -125 209 -119
rect 175 -187 209 -163
rect 175 -197 209 -187
rect 175 -255 209 -235
rect 175 -269 209 -255
rect 271 255 305 269
rect 271 235 305 255
rect 271 187 305 197
rect 271 163 305 187
rect 271 119 305 125
rect 271 91 305 119
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect 271 -119 305 -91
rect 271 -125 305 -119
rect 271 -187 305 -163
rect 271 -197 305 -187
rect 271 -255 305 -235
rect 271 -269 305 -255
rect 367 255 401 269
rect 367 235 401 255
rect 367 187 401 197
rect 367 163 401 187
rect 367 119 401 125
rect 367 91 401 119
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 367 -119 401 -91
rect 367 -125 401 -119
rect 367 -187 401 -163
rect 367 -197 401 -187
rect 367 -255 401 -235
rect 367 -269 401 -255
rect 463 255 497 269
rect 463 235 497 255
rect 463 187 497 197
rect 463 163 497 187
rect 463 119 497 125
rect 463 91 497 119
rect 463 51 497 53
rect 463 19 497 51
rect 463 -51 497 -19
rect 463 -53 497 -51
rect 463 -119 497 -91
rect 463 -125 497 -119
rect 463 -187 497 -163
rect 463 -197 497 -187
rect 463 -255 497 -235
rect 463 -269 497 -255
rect 559 255 593 269
rect 559 235 593 255
rect 559 187 593 197
rect 559 163 593 187
rect 559 119 593 125
rect 559 91 593 119
rect 559 51 593 53
rect 559 19 593 51
rect 559 -51 593 -19
rect 559 -53 593 -51
rect 559 -119 593 -91
rect 559 -125 593 -119
rect 559 -187 593 -163
rect 559 -197 593 -187
rect 559 -255 593 -235
rect 559 -269 593 -255
rect 655 255 689 269
rect 655 235 689 255
rect 655 187 689 197
rect 655 163 689 187
rect 655 119 689 125
rect 655 91 689 119
rect 655 51 689 53
rect 655 19 689 51
rect 655 -51 689 -19
rect 655 -53 689 -51
rect 655 -119 689 -91
rect 655 -125 689 -119
rect 655 -187 689 -163
rect 655 -197 689 -187
rect 655 -255 689 -235
rect 655 -269 689 -255
rect 751 255 785 269
rect 751 235 785 255
rect 751 187 785 197
rect 751 163 785 187
rect 751 119 785 125
rect 751 91 785 119
rect 751 51 785 53
rect 751 19 785 51
rect 751 -51 785 -19
rect 751 -53 785 -51
rect 751 -119 785 -91
rect 751 -125 785 -119
rect 751 -187 785 -163
rect 751 -197 785 -187
rect 751 -255 785 -235
rect 751 -269 785 -255
rect 847 255 881 269
rect 847 235 881 255
rect 847 187 881 197
rect 847 163 881 187
rect 847 119 881 125
rect 847 91 881 119
rect 847 51 881 53
rect 847 19 881 51
rect 847 -51 881 -19
rect 847 -53 881 -51
rect 847 -119 881 -91
rect 847 -125 881 -119
rect 847 -187 881 -163
rect 847 -197 881 -187
rect 847 -255 881 -235
rect 847 -269 881 -255
rect 943 255 977 269
rect 943 235 977 255
rect 943 187 977 197
rect 943 163 977 187
rect 943 119 977 125
rect 943 91 977 119
rect 943 51 977 53
rect 943 19 977 51
rect 943 -51 977 -19
rect 943 -53 977 -51
rect 943 -119 977 -91
rect 943 -125 977 -119
rect 943 -187 977 -163
rect 943 -197 977 -187
rect 943 -255 977 -235
rect 943 -269 977 -255
rect 1039 255 1073 269
rect 1039 235 1073 255
rect 1039 187 1073 197
rect 1039 163 1073 187
rect 1039 119 1073 125
rect 1039 91 1073 119
rect 1039 51 1073 53
rect 1039 19 1073 51
rect 1039 -51 1073 -19
rect 1039 -53 1073 -51
rect 1039 -119 1073 -91
rect 1039 -125 1073 -119
rect 1039 -187 1073 -163
rect 1039 -197 1073 -187
rect 1039 -255 1073 -235
rect 1039 -269 1073 -255
rect 1135 255 1169 269
rect 1135 235 1169 255
rect 1135 187 1169 197
rect 1135 163 1169 187
rect 1135 119 1169 125
rect 1135 91 1169 119
rect 1135 51 1169 53
rect 1135 19 1169 51
rect 1135 -51 1169 -19
rect 1135 -53 1169 -51
rect 1135 -119 1169 -91
rect 1135 -125 1169 -119
rect 1135 -187 1169 -163
rect 1135 -197 1169 -187
rect 1135 -255 1169 -235
rect 1135 -269 1169 -255
rect 1231 255 1265 269
rect 1231 235 1265 255
rect 1231 187 1265 197
rect 1231 163 1265 187
rect 1231 119 1265 125
rect 1231 91 1265 119
rect 1231 51 1265 53
rect 1231 19 1265 51
rect 1231 -51 1265 -19
rect 1231 -53 1265 -51
rect 1231 -119 1265 -91
rect 1231 -125 1265 -119
rect 1231 -187 1265 -163
rect 1231 -197 1265 -187
rect 1231 -255 1265 -235
rect 1231 -269 1265 -255
rect 1327 255 1361 269
rect 1327 235 1361 255
rect 1327 187 1361 197
rect 1327 163 1361 187
rect 1327 119 1361 125
rect 1327 91 1361 119
rect 1327 51 1361 53
rect 1327 19 1361 51
rect 1327 -51 1361 -19
rect 1327 -53 1361 -51
rect 1327 -119 1361 -91
rect 1327 -125 1361 -119
rect 1327 -187 1361 -163
rect 1327 -197 1361 -187
rect 1327 -255 1361 -235
rect 1327 -269 1361 -255
rect 1423 255 1457 269
rect 1423 235 1457 255
rect 1423 187 1457 197
rect 1423 163 1457 187
rect 1423 119 1457 125
rect 1423 91 1457 119
rect 1423 51 1457 53
rect 1423 19 1457 51
rect 1423 -51 1457 -19
rect 1423 -53 1457 -51
rect 1423 -119 1457 -91
rect 1423 -125 1457 -119
rect 1423 -187 1457 -163
rect 1423 -197 1457 -187
rect 1423 -255 1457 -235
rect 1423 -269 1457 -255
rect 1519 255 1553 269
rect 1519 235 1553 255
rect 1519 187 1553 197
rect 1519 163 1553 187
rect 1519 119 1553 125
rect 1519 91 1553 119
rect 1519 51 1553 53
rect 1519 19 1553 51
rect 1519 -51 1553 -19
rect 1519 -53 1553 -51
rect 1519 -119 1553 -91
rect 1519 -125 1553 -119
rect 1519 -187 1553 -163
rect 1519 -197 1553 -187
rect 1519 -255 1553 -235
rect 1519 -269 1553 -255
rect 1615 255 1649 269
rect 1615 235 1649 255
rect 1615 187 1649 197
rect 1615 163 1649 187
rect 1615 119 1649 125
rect 1615 91 1649 119
rect 1615 51 1649 53
rect 1615 19 1649 51
rect 1615 -51 1649 -19
rect 1615 -53 1649 -51
rect 1615 -119 1649 -91
rect 1615 -125 1649 -119
rect 1615 -187 1649 -163
rect 1615 -197 1649 -187
rect 1615 -255 1649 -235
rect 1615 -269 1649 -255
rect 1711 255 1745 269
rect 1711 235 1745 255
rect 1711 187 1745 197
rect 1711 163 1745 187
rect 1711 119 1745 125
rect 1711 91 1745 119
rect 1711 51 1745 53
rect 1711 19 1745 51
rect 1711 -51 1745 -19
rect 1711 -53 1745 -51
rect 1711 -119 1745 -91
rect 1711 -125 1745 -119
rect 1711 -187 1745 -163
rect 1711 -197 1745 -187
rect 1711 -255 1745 -235
rect 1711 -269 1745 -255
rect 1807 255 1841 269
rect 1807 235 1841 255
rect 1807 187 1841 197
rect 1807 163 1841 187
rect 1807 119 1841 125
rect 1807 91 1841 119
rect 1807 51 1841 53
rect 1807 19 1841 51
rect 1807 -51 1841 -19
rect 1807 -53 1841 -51
rect 1807 -119 1841 -91
rect 1807 -125 1841 -119
rect 1807 -187 1841 -163
rect 1807 -197 1841 -187
rect 1807 -255 1841 -235
rect 1807 -269 1841 -255
rect 1903 255 1937 269
rect 1903 235 1937 255
rect 1903 187 1937 197
rect 1903 163 1937 187
rect 1903 119 1937 125
rect 1903 91 1937 119
rect 1903 51 1937 53
rect 1903 19 1937 51
rect 1903 -51 1937 -19
rect 1903 -53 1937 -51
rect 1903 -119 1937 -91
rect 1903 -125 1937 -119
rect 1903 -187 1937 -163
rect 1903 -197 1937 -187
rect 1903 -255 1937 -235
rect 1903 -269 1937 -255
rect 1999 255 2033 269
rect 1999 235 2033 255
rect 1999 187 2033 197
rect 1999 163 2033 187
rect 1999 119 2033 125
rect 1999 91 2033 119
rect 1999 51 2033 53
rect 1999 19 2033 51
rect 1999 -51 2033 -19
rect 1999 -53 2033 -51
rect 1999 -119 2033 -91
rect 1999 -125 2033 -119
rect 1999 -187 2033 -163
rect 1999 -197 2033 -187
rect 1999 -255 2033 -235
rect 1999 -269 2033 -255
rect -1985 -372 -1951 -338
rect -1793 -372 -1759 -338
rect -1601 -372 -1567 -338
rect -1409 -372 -1375 -338
rect -1217 -372 -1183 -338
rect -1025 -372 -991 -338
rect -833 -372 -799 -338
rect -641 -372 -607 -338
rect -449 -372 -415 -338
rect -257 -372 -223 -338
rect -65 -372 -31 -338
rect 127 -372 161 -338
rect 319 -372 353 -338
rect 511 -372 545 -338
rect 703 -372 737 -338
rect 895 -372 929 -338
rect 1087 -372 1121 -338
rect 1279 -372 1313 -338
rect 1471 -372 1505 -338
rect 1663 -372 1697 -338
rect 1855 -372 1889 -338
<< metal1 >>
rect -1901 372 -1843 378
rect -1901 338 -1889 372
rect -1855 338 -1843 372
rect -1901 332 -1843 338
rect -1709 372 -1651 378
rect -1709 338 -1697 372
rect -1663 338 -1651 372
rect -1709 332 -1651 338
rect -1517 372 -1459 378
rect -1517 338 -1505 372
rect -1471 338 -1459 372
rect -1517 332 -1459 338
rect -1325 372 -1267 378
rect -1325 338 -1313 372
rect -1279 338 -1267 372
rect -1325 332 -1267 338
rect -1133 372 -1075 378
rect -1133 338 -1121 372
rect -1087 338 -1075 372
rect -1133 332 -1075 338
rect -941 372 -883 378
rect -941 338 -929 372
rect -895 338 -883 372
rect -941 332 -883 338
rect -749 372 -691 378
rect -749 338 -737 372
rect -703 338 -691 372
rect -749 332 -691 338
rect -557 372 -499 378
rect -557 338 -545 372
rect -511 338 -499 372
rect -557 332 -499 338
rect -365 372 -307 378
rect -365 338 -353 372
rect -319 338 -307 372
rect -365 332 -307 338
rect -173 372 -115 378
rect -173 338 -161 372
rect -127 338 -115 372
rect -173 332 -115 338
rect 19 372 77 378
rect 19 338 31 372
rect 65 338 77 372
rect 19 332 77 338
rect 211 372 269 378
rect 211 338 223 372
rect 257 338 269 372
rect 211 332 269 338
rect 403 372 461 378
rect 403 338 415 372
rect 449 338 461 372
rect 403 332 461 338
rect 595 372 653 378
rect 595 338 607 372
rect 641 338 653 372
rect 595 332 653 338
rect 787 372 845 378
rect 787 338 799 372
rect 833 338 845 372
rect 787 332 845 338
rect 979 372 1037 378
rect 979 338 991 372
rect 1025 338 1037 372
rect 979 332 1037 338
rect 1171 372 1229 378
rect 1171 338 1183 372
rect 1217 338 1229 372
rect 1171 332 1229 338
rect 1363 372 1421 378
rect 1363 338 1375 372
rect 1409 338 1421 372
rect 1363 332 1421 338
rect 1555 372 1613 378
rect 1555 338 1567 372
rect 1601 338 1613 372
rect 1555 332 1613 338
rect 1747 372 1805 378
rect 1747 338 1759 372
rect 1793 338 1805 372
rect 1747 332 1805 338
rect 1939 372 1997 378
rect 1939 338 1951 372
rect 1985 338 1997 372
rect 1939 332 1997 338
rect -2039 269 -1993 300
rect -2039 235 -2033 269
rect -1999 235 -1993 269
rect -2039 197 -1993 235
rect -2039 163 -2033 197
rect -1999 163 -1993 197
rect -2039 125 -1993 163
rect -2039 91 -2033 125
rect -1999 91 -1993 125
rect -2039 53 -1993 91
rect -2039 19 -2033 53
rect -1999 19 -1993 53
rect -2039 -19 -1993 19
rect -2039 -53 -2033 -19
rect -1999 -53 -1993 -19
rect -2039 -91 -1993 -53
rect -2039 -125 -2033 -91
rect -1999 -125 -1993 -91
rect -2039 -163 -1993 -125
rect -2039 -197 -2033 -163
rect -1999 -197 -1993 -163
rect -2039 -235 -1993 -197
rect -2039 -269 -2033 -235
rect -1999 -269 -1993 -235
rect -2039 -300 -1993 -269
rect -1943 269 -1897 300
rect -1943 235 -1937 269
rect -1903 235 -1897 269
rect -1943 197 -1897 235
rect -1943 163 -1937 197
rect -1903 163 -1897 197
rect -1943 125 -1897 163
rect -1943 91 -1937 125
rect -1903 91 -1897 125
rect -1943 53 -1897 91
rect -1943 19 -1937 53
rect -1903 19 -1897 53
rect -1943 -19 -1897 19
rect -1943 -53 -1937 -19
rect -1903 -53 -1897 -19
rect -1943 -91 -1897 -53
rect -1943 -125 -1937 -91
rect -1903 -125 -1897 -91
rect -1943 -163 -1897 -125
rect -1943 -197 -1937 -163
rect -1903 -197 -1897 -163
rect -1943 -235 -1897 -197
rect -1943 -269 -1937 -235
rect -1903 -269 -1897 -235
rect -1943 -300 -1897 -269
rect -1847 269 -1801 300
rect -1847 235 -1841 269
rect -1807 235 -1801 269
rect -1847 197 -1801 235
rect -1847 163 -1841 197
rect -1807 163 -1801 197
rect -1847 125 -1801 163
rect -1847 91 -1841 125
rect -1807 91 -1801 125
rect -1847 53 -1801 91
rect -1847 19 -1841 53
rect -1807 19 -1801 53
rect -1847 -19 -1801 19
rect -1847 -53 -1841 -19
rect -1807 -53 -1801 -19
rect -1847 -91 -1801 -53
rect -1847 -125 -1841 -91
rect -1807 -125 -1801 -91
rect -1847 -163 -1801 -125
rect -1847 -197 -1841 -163
rect -1807 -197 -1801 -163
rect -1847 -235 -1801 -197
rect -1847 -269 -1841 -235
rect -1807 -269 -1801 -235
rect -1847 -300 -1801 -269
rect -1751 269 -1705 300
rect -1751 235 -1745 269
rect -1711 235 -1705 269
rect -1751 197 -1705 235
rect -1751 163 -1745 197
rect -1711 163 -1705 197
rect -1751 125 -1705 163
rect -1751 91 -1745 125
rect -1711 91 -1705 125
rect -1751 53 -1705 91
rect -1751 19 -1745 53
rect -1711 19 -1705 53
rect -1751 -19 -1705 19
rect -1751 -53 -1745 -19
rect -1711 -53 -1705 -19
rect -1751 -91 -1705 -53
rect -1751 -125 -1745 -91
rect -1711 -125 -1705 -91
rect -1751 -163 -1705 -125
rect -1751 -197 -1745 -163
rect -1711 -197 -1705 -163
rect -1751 -235 -1705 -197
rect -1751 -269 -1745 -235
rect -1711 -269 -1705 -235
rect -1751 -300 -1705 -269
rect -1655 269 -1609 300
rect -1655 235 -1649 269
rect -1615 235 -1609 269
rect -1655 197 -1609 235
rect -1655 163 -1649 197
rect -1615 163 -1609 197
rect -1655 125 -1609 163
rect -1655 91 -1649 125
rect -1615 91 -1609 125
rect -1655 53 -1609 91
rect -1655 19 -1649 53
rect -1615 19 -1609 53
rect -1655 -19 -1609 19
rect -1655 -53 -1649 -19
rect -1615 -53 -1609 -19
rect -1655 -91 -1609 -53
rect -1655 -125 -1649 -91
rect -1615 -125 -1609 -91
rect -1655 -163 -1609 -125
rect -1655 -197 -1649 -163
rect -1615 -197 -1609 -163
rect -1655 -235 -1609 -197
rect -1655 -269 -1649 -235
rect -1615 -269 -1609 -235
rect -1655 -300 -1609 -269
rect -1559 269 -1513 300
rect -1559 235 -1553 269
rect -1519 235 -1513 269
rect -1559 197 -1513 235
rect -1559 163 -1553 197
rect -1519 163 -1513 197
rect -1559 125 -1513 163
rect -1559 91 -1553 125
rect -1519 91 -1513 125
rect -1559 53 -1513 91
rect -1559 19 -1553 53
rect -1519 19 -1513 53
rect -1559 -19 -1513 19
rect -1559 -53 -1553 -19
rect -1519 -53 -1513 -19
rect -1559 -91 -1513 -53
rect -1559 -125 -1553 -91
rect -1519 -125 -1513 -91
rect -1559 -163 -1513 -125
rect -1559 -197 -1553 -163
rect -1519 -197 -1513 -163
rect -1559 -235 -1513 -197
rect -1559 -269 -1553 -235
rect -1519 -269 -1513 -235
rect -1559 -300 -1513 -269
rect -1463 269 -1417 300
rect -1463 235 -1457 269
rect -1423 235 -1417 269
rect -1463 197 -1417 235
rect -1463 163 -1457 197
rect -1423 163 -1417 197
rect -1463 125 -1417 163
rect -1463 91 -1457 125
rect -1423 91 -1417 125
rect -1463 53 -1417 91
rect -1463 19 -1457 53
rect -1423 19 -1417 53
rect -1463 -19 -1417 19
rect -1463 -53 -1457 -19
rect -1423 -53 -1417 -19
rect -1463 -91 -1417 -53
rect -1463 -125 -1457 -91
rect -1423 -125 -1417 -91
rect -1463 -163 -1417 -125
rect -1463 -197 -1457 -163
rect -1423 -197 -1417 -163
rect -1463 -235 -1417 -197
rect -1463 -269 -1457 -235
rect -1423 -269 -1417 -235
rect -1463 -300 -1417 -269
rect -1367 269 -1321 300
rect -1367 235 -1361 269
rect -1327 235 -1321 269
rect -1367 197 -1321 235
rect -1367 163 -1361 197
rect -1327 163 -1321 197
rect -1367 125 -1321 163
rect -1367 91 -1361 125
rect -1327 91 -1321 125
rect -1367 53 -1321 91
rect -1367 19 -1361 53
rect -1327 19 -1321 53
rect -1367 -19 -1321 19
rect -1367 -53 -1361 -19
rect -1327 -53 -1321 -19
rect -1367 -91 -1321 -53
rect -1367 -125 -1361 -91
rect -1327 -125 -1321 -91
rect -1367 -163 -1321 -125
rect -1367 -197 -1361 -163
rect -1327 -197 -1321 -163
rect -1367 -235 -1321 -197
rect -1367 -269 -1361 -235
rect -1327 -269 -1321 -235
rect -1367 -300 -1321 -269
rect -1271 269 -1225 300
rect -1271 235 -1265 269
rect -1231 235 -1225 269
rect -1271 197 -1225 235
rect -1271 163 -1265 197
rect -1231 163 -1225 197
rect -1271 125 -1225 163
rect -1271 91 -1265 125
rect -1231 91 -1225 125
rect -1271 53 -1225 91
rect -1271 19 -1265 53
rect -1231 19 -1225 53
rect -1271 -19 -1225 19
rect -1271 -53 -1265 -19
rect -1231 -53 -1225 -19
rect -1271 -91 -1225 -53
rect -1271 -125 -1265 -91
rect -1231 -125 -1225 -91
rect -1271 -163 -1225 -125
rect -1271 -197 -1265 -163
rect -1231 -197 -1225 -163
rect -1271 -235 -1225 -197
rect -1271 -269 -1265 -235
rect -1231 -269 -1225 -235
rect -1271 -300 -1225 -269
rect -1175 269 -1129 300
rect -1175 235 -1169 269
rect -1135 235 -1129 269
rect -1175 197 -1129 235
rect -1175 163 -1169 197
rect -1135 163 -1129 197
rect -1175 125 -1129 163
rect -1175 91 -1169 125
rect -1135 91 -1129 125
rect -1175 53 -1129 91
rect -1175 19 -1169 53
rect -1135 19 -1129 53
rect -1175 -19 -1129 19
rect -1175 -53 -1169 -19
rect -1135 -53 -1129 -19
rect -1175 -91 -1129 -53
rect -1175 -125 -1169 -91
rect -1135 -125 -1129 -91
rect -1175 -163 -1129 -125
rect -1175 -197 -1169 -163
rect -1135 -197 -1129 -163
rect -1175 -235 -1129 -197
rect -1175 -269 -1169 -235
rect -1135 -269 -1129 -235
rect -1175 -300 -1129 -269
rect -1079 269 -1033 300
rect -1079 235 -1073 269
rect -1039 235 -1033 269
rect -1079 197 -1033 235
rect -1079 163 -1073 197
rect -1039 163 -1033 197
rect -1079 125 -1033 163
rect -1079 91 -1073 125
rect -1039 91 -1033 125
rect -1079 53 -1033 91
rect -1079 19 -1073 53
rect -1039 19 -1033 53
rect -1079 -19 -1033 19
rect -1079 -53 -1073 -19
rect -1039 -53 -1033 -19
rect -1079 -91 -1033 -53
rect -1079 -125 -1073 -91
rect -1039 -125 -1033 -91
rect -1079 -163 -1033 -125
rect -1079 -197 -1073 -163
rect -1039 -197 -1033 -163
rect -1079 -235 -1033 -197
rect -1079 -269 -1073 -235
rect -1039 -269 -1033 -235
rect -1079 -300 -1033 -269
rect -983 269 -937 300
rect -983 235 -977 269
rect -943 235 -937 269
rect -983 197 -937 235
rect -983 163 -977 197
rect -943 163 -937 197
rect -983 125 -937 163
rect -983 91 -977 125
rect -943 91 -937 125
rect -983 53 -937 91
rect -983 19 -977 53
rect -943 19 -937 53
rect -983 -19 -937 19
rect -983 -53 -977 -19
rect -943 -53 -937 -19
rect -983 -91 -937 -53
rect -983 -125 -977 -91
rect -943 -125 -937 -91
rect -983 -163 -937 -125
rect -983 -197 -977 -163
rect -943 -197 -937 -163
rect -983 -235 -937 -197
rect -983 -269 -977 -235
rect -943 -269 -937 -235
rect -983 -300 -937 -269
rect -887 269 -841 300
rect -887 235 -881 269
rect -847 235 -841 269
rect -887 197 -841 235
rect -887 163 -881 197
rect -847 163 -841 197
rect -887 125 -841 163
rect -887 91 -881 125
rect -847 91 -841 125
rect -887 53 -841 91
rect -887 19 -881 53
rect -847 19 -841 53
rect -887 -19 -841 19
rect -887 -53 -881 -19
rect -847 -53 -841 -19
rect -887 -91 -841 -53
rect -887 -125 -881 -91
rect -847 -125 -841 -91
rect -887 -163 -841 -125
rect -887 -197 -881 -163
rect -847 -197 -841 -163
rect -887 -235 -841 -197
rect -887 -269 -881 -235
rect -847 -269 -841 -235
rect -887 -300 -841 -269
rect -791 269 -745 300
rect -791 235 -785 269
rect -751 235 -745 269
rect -791 197 -745 235
rect -791 163 -785 197
rect -751 163 -745 197
rect -791 125 -745 163
rect -791 91 -785 125
rect -751 91 -745 125
rect -791 53 -745 91
rect -791 19 -785 53
rect -751 19 -745 53
rect -791 -19 -745 19
rect -791 -53 -785 -19
rect -751 -53 -745 -19
rect -791 -91 -745 -53
rect -791 -125 -785 -91
rect -751 -125 -745 -91
rect -791 -163 -745 -125
rect -791 -197 -785 -163
rect -751 -197 -745 -163
rect -791 -235 -745 -197
rect -791 -269 -785 -235
rect -751 -269 -745 -235
rect -791 -300 -745 -269
rect -695 269 -649 300
rect -695 235 -689 269
rect -655 235 -649 269
rect -695 197 -649 235
rect -695 163 -689 197
rect -655 163 -649 197
rect -695 125 -649 163
rect -695 91 -689 125
rect -655 91 -649 125
rect -695 53 -649 91
rect -695 19 -689 53
rect -655 19 -649 53
rect -695 -19 -649 19
rect -695 -53 -689 -19
rect -655 -53 -649 -19
rect -695 -91 -649 -53
rect -695 -125 -689 -91
rect -655 -125 -649 -91
rect -695 -163 -649 -125
rect -695 -197 -689 -163
rect -655 -197 -649 -163
rect -695 -235 -649 -197
rect -695 -269 -689 -235
rect -655 -269 -649 -235
rect -695 -300 -649 -269
rect -599 269 -553 300
rect -599 235 -593 269
rect -559 235 -553 269
rect -599 197 -553 235
rect -599 163 -593 197
rect -559 163 -553 197
rect -599 125 -553 163
rect -599 91 -593 125
rect -559 91 -553 125
rect -599 53 -553 91
rect -599 19 -593 53
rect -559 19 -553 53
rect -599 -19 -553 19
rect -599 -53 -593 -19
rect -559 -53 -553 -19
rect -599 -91 -553 -53
rect -599 -125 -593 -91
rect -559 -125 -553 -91
rect -599 -163 -553 -125
rect -599 -197 -593 -163
rect -559 -197 -553 -163
rect -599 -235 -553 -197
rect -599 -269 -593 -235
rect -559 -269 -553 -235
rect -599 -300 -553 -269
rect -503 269 -457 300
rect -503 235 -497 269
rect -463 235 -457 269
rect -503 197 -457 235
rect -503 163 -497 197
rect -463 163 -457 197
rect -503 125 -457 163
rect -503 91 -497 125
rect -463 91 -457 125
rect -503 53 -457 91
rect -503 19 -497 53
rect -463 19 -457 53
rect -503 -19 -457 19
rect -503 -53 -497 -19
rect -463 -53 -457 -19
rect -503 -91 -457 -53
rect -503 -125 -497 -91
rect -463 -125 -457 -91
rect -503 -163 -457 -125
rect -503 -197 -497 -163
rect -463 -197 -457 -163
rect -503 -235 -457 -197
rect -503 -269 -497 -235
rect -463 -269 -457 -235
rect -503 -300 -457 -269
rect -407 269 -361 300
rect -407 235 -401 269
rect -367 235 -361 269
rect -407 197 -361 235
rect -407 163 -401 197
rect -367 163 -361 197
rect -407 125 -361 163
rect -407 91 -401 125
rect -367 91 -361 125
rect -407 53 -361 91
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -91 -361 -53
rect -407 -125 -401 -91
rect -367 -125 -361 -91
rect -407 -163 -361 -125
rect -407 -197 -401 -163
rect -367 -197 -361 -163
rect -407 -235 -361 -197
rect -407 -269 -401 -235
rect -367 -269 -361 -235
rect -407 -300 -361 -269
rect -311 269 -265 300
rect -311 235 -305 269
rect -271 235 -265 269
rect -311 197 -265 235
rect -311 163 -305 197
rect -271 163 -265 197
rect -311 125 -265 163
rect -311 91 -305 125
rect -271 91 -265 125
rect -311 53 -265 91
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -91 -265 -53
rect -311 -125 -305 -91
rect -271 -125 -265 -91
rect -311 -163 -265 -125
rect -311 -197 -305 -163
rect -271 -197 -265 -163
rect -311 -235 -265 -197
rect -311 -269 -305 -235
rect -271 -269 -265 -235
rect -311 -300 -265 -269
rect -215 269 -169 300
rect -215 235 -209 269
rect -175 235 -169 269
rect -215 197 -169 235
rect -215 163 -209 197
rect -175 163 -169 197
rect -215 125 -169 163
rect -215 91 -209 125
rect -175 91 -169 125
rect -215 53 -169 91
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -91 -169 -53
rect -215 -125 -209 -91
rect -175 -125 -169 -91
rect -215 -163 -169 -125
rect -215 -197 -209 -163
rect -175 -197 -169 -163
rect -215 -235 -169 -197
rect -215 -269 -209 -235
rect -175 -269 -169 -235
rect -215 -300 -169 -269
rect -119 269 -73 300
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -300 -73 -269
rect -23 269 23 300
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -300 23 -269
rect 73 269 119 300
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -300 119 -269
rect 169 269 215 300
rect 169 235 175 269
rect 209 235 215 269
rect 169 197 215 235
rect 169 163 175 197
rect 209 163 215 197
rect 169 125 215 163
rect 169 91 175 125
rect 209 91 215 125
rect 169 53 215 91
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -91 215 -53
rect 169 -125 175 -91
rect 209 -125 215 -91
rect 169 -163 215 -125
rect 169 -197 175 -163
rect 209 -197 215 -163
rect 169 -235 215 -197
rect 169 -269 175 -235
rect 209 -269 215 -235
rect 169 -300 215 -269
rect 265 269 311 300
rect 265 235 271 269
rect 305 235 311 269
rect 265 197 311 235
rect 265 163 271 197
rect 305 163 311 197
rect 265 125 311 163
rect 265 91 271 125
rect 305 91 311 125
rect 265 53 311 91
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -91 311 -53
rect 265 -125 271 -91
rect 305 -125 311 -91
rect 265 -163 311 -125
rect 265 -197 271 -163
rect 305 -197 311 -163
rect 265 -235 311 -197
rect 265 -269 271 -235
rect 305 -269 311 -235
rect 265 -300 311 -269
rect 361 269 407 300
rect 361 235 367 269
rect 401 235 407 269
rect 361 197 407 235
rect 361 163 367 197
rect 401 163 407 197
rect 361 125 407 163
rect 361 91 367 125
rect 401 91 407 125
rect 361 53 407 91
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -91 407 -53
rect 361 -125 367 -91
rect 401 -125 407 -91
rect 361 -163 407 -125
rect 361 -197 367 -163
rect 401 -197 407 -163
rect 361 -235 407 -197
rect 361 -269 367 -235
rect 401 -269 407 -235
rect 361 -300 407 -269
rect 457 269 503 300
rect 457 235 463 269
rect 497 235 503 269
rect 457 197 503 235
rect 457 163 463 197
rect 497 163 503 197
rect 457 125 503 163
rect 457 91 463 125
rect 497 91 503 125
rect 457 53 503 91
rect 457 19 463 53
rect 497 19 503 53
rect 457 -19 503 19
rect 457 -53 463 -19
rect 497 -53 503 -19
rect 457 -91 503 -53
rect 457 -125 463 -91
rect 497 -125 503 -91
rect 457 -163 503 -125
rect 457 -197 463 -163
rect 497 -197 503 -163
rect 457 -235 503 -197
rect 457 -269 463 -235
rect 497 -269 503 -235
rect 457 -300 503 -269
rect 553 269 599 300
rect 553 235 559 269
rect 593 235 599 269
rect 553 197 599 235
rect 553 163 559 197
rect 593 163 599 197
rect 553 125 599 163
rect 553 91 559 125
rect 593 91 599 125
rect 553 53 599 91
rect 553 19 559 53
rect 593 19 599 53
rect 553 -19 599 19
rect 553 -53 559 -19
rect 593 -53 599 -19
rect 553 -91 599 -53
rect 553 -125 559 -91
rect 593 -125 599 -91
rect 553 -163 599 -125
rect 553 -197 559 -163
rect 593 -197 599 -163
rect 553 -235 599 -197
rect 553 -269 559 -235
rect 593 -269 599 -235
rect 553 -300 599 -269
rect 649 269 695 300
rect 649 235 655 269
rect 689 235 695 269
rect 649 197 695 235
rect 649 163 655 197
rect 689 163 695 197
rect 649 125 695 163
rect 649 91 655 125
rect 689 91 695 125
rect 649 53 695 91
rect 649 19 655 53
rect 689 19 695 53
rect 649 -19 695 19
rect 649 -53 655 -19
rect 689 -53 695 -19
rect 649 -91 695 -53
rect 649 -125 655 -91
rect 689 -125 695 -91
rect 649 -163 695 -125
rect 649 -197 655 -163
rect 689 -197 695 -163
rect 649 -235 695 -197
rect 649 -269 655 -235
rect 689 -269 695 -235
rect 649 -300 695 -269
rect 745 269 791 300
rect 745 235 751 269
rect 785 235 791 269
rect 745 197 791 235
rect 745 163 751 197
rect 785 163 791 197
rect 745 125 791 163
rect 745 91 751 125
rect 785 91 791 125
rect 745 53 791 91
rect 745 19 751 53
rect 785 19 791 53
rect 745 -19 791 19
rect 745 -53 751 -19
rect 785 -53 791 -19
rect 745 -91 791 -53
rect 745 -125 751 -91
rect 785 -125 791 -91
rect 745 -163 791 -125
rect 745 -197 751 -163
rect 785 -197 791 -163
rect 745 -235 791 -197
rect 745 -269 751 -235
rect 785 -269 791 -235
rect 745 -300 791 -269
rect 841 269 887 300
rect 841 235 847 269
rect 881 235 887 269
rect 841 197 887 235
rect 841 163 847 197
rect 881 163 887 197
rect 841 125 887 163
rect 841 91 847 125
rect 881 91 887 125
rect 841 53 887 91
rect 841 19 847 53
rect 881 19 887 53
rect 841 -19 887 19
rect 841 -53 847 -19
rect 881 -53 887 -19
rect 841 -91 887 -53
rect 841 -125 847 -91
rect 881 -125 887 -91
rect 841 -163 887 -125
rect 841 -197 847 -163
rect 881 -197 887 -163
rect 841 -235 887 -197
rect 841 -269 847 -235
rect 881 -269 887 -235
rect 841 -300 887 -269
rect 937 269 983 300
rect 937 235 943 269
rect 977 235 983 269
rect 937 197 983 235
rect 937 163 943 197
rect 977 163 983 197
rect 937 125 983 163
rect 937 91 943 125
rect 977 91 983 125
rect 937 53 983 91
rect 937 19 943 53
rect 977 19 983 53
rect 937 -19 983 19
rect 937 -53 943 -19
rect 977 -53 983 -19
rect 937 -91 983 -53
rect 937 -125 943 -91
rect 977 -125 983 -91
rect 937 -163 983 -125
rect 937 -197 943 -163
rect 977 -197 983 -163
rect 937 -235 983 -197
rect 937 -269 943 -235
rect 977 -269 983 -235
rect 937 -300 983 -269
rect 1033 269 1079 300
rect 1033 235 1039 269
rect 1073 235 1079 269
rect 1033 197 1079 235
rect 1033 163 1039 197
rect 1073 163 1079 197
rect 1033 125 1079 163
rect 1033 91 1039 125
rect 1073 91 1079 125
rect 1033 53 1079 91
rect 1033 19 1039 53
rect 1073 19 1079 53
rect 1033 -19 1079 19
rect 1033 -53 1039 -19
rect 1073 -53 1079 -19
rect 1033 -91 1079 -53
rect 1033 -125 1039 -91
rect 1073 -125 1079 -91
rect 1033 -163 1079 -125
rect 1033 -197 1039 -163
rect 1073 -197 1079 -163
rect 1033 -235 1079 -197
rect 1033 -269 1039 -235
rect 1073 -269 1079 -235
rect 1033 -300 1079 -269
rect 1129 269 1175 300
rect 1129 235 1135 269
rect 1169 235 1175 269
rect 1129 197 1175 235
rect 1129 163 1135 197
rect 1169 163 1175 197
rect 1129 125 1175 163
rect 1129 91 1135 125
rect 1169 91 1175 125
rect 1129 53 1175 91
rect 1129 19 1135 53
rect 1169 19 1175 53
rect 1129 -19 1175 19
rect 1129 -53 1135 -19
rect 1169 -53 1175 -19
rect 1129 -91 1175 -53
rect 1129 -125 1135 -91
rect 1169 -125 1175 -91
rect 1129 -163 1175 -125
rect 1129 -197 1135 -163
rect 1169 -197 1175 -163
rect 1129 -235 1175 -197
rect 1129 -269 1135 -235
rect 1169 -269 1175 -235
rect 1129 -300 1175 -269
rect 1225 269 1271 300
rect 1225 235 1231 269
rect 1265 235 1271 269
rect 1225 197 1271 235
rect 1225 163 1231 197
rect 1265 163 1271 197
rect 1225 125 1271 163
rect 1225 91 1231 125
rect 1265 91 1271 125
rect 1225 53 1271 91
rect 1225 19 1231 53
rect 1265 19 1271 53
rect 1225 -19 1271 19
rect 1225 -53 1231 -19
rect 1265 -53 1271 -19
rect 1225 -91 1271 -53
rect 1225 -125 1231 -91
rect 1265 -125 1271 -91
rect 1225 -163 1271 -125
rect 1225 -197 1231 -163
rect 1265 -197 1271 -163
rect 1225 -235 1271 -197
rect 1225 -269 1231 -235
rect 1265 -269 1271 -235
rect 1225 -300 1271 -269
rect 1321 269 1367 300
rect 1321 235 1327 269
rect 1361 235 1367 269
rect 1321 197 1367 235
rect 1321 163 1327 197
rect 1361 163 1367 197
rect 1321 125 1367 163
rect 1321 91 1327 125
rect 1361 91 1367 125
rect 1321 53 1367 91
rect 1321 19 1327 53
rect 1361 19 1367 53
rect 1321 -19 1367 19
rect 1321 -53 1327 -19
rect 1361 -53 1367 -19
rect 1321 -91 1367 -53
rect 1321 -125 1327 -91
rect 1361 -125 1367 -91
rect 1321 -163 1367 -125
rect 1321 -197 1327 -163
rect 1361 -197 1367 -163
rect 1321 -235 1367 -197
rect 1321 -269 1327 -235
rect 1361 -269 1367 -235
rect 1321 -300 1367 -269
rect 1417 269 1463 300
rect 1417 235 1423 269
rect 1457 235 1463 269
rect 1417 197 1463 235
rect 1417 163 1423 197
rect 1457 163 1463 197
rect 1417 125 1463 163
rect 1417 91 1423 125
rect 1457 91 1463 125
rect 1417 53 1463 91
rect 1417 19 1423 53
rect 1457 19 1463 53
rect 1417 -19 1463 19
rect 1417 -53 1423 -19
rect 1457 -53 1463 -19
rect 1417 -91 1463 -53
rect 1417 -125 1423 -91
rect 1457 -125 1463 -91
rect 1417 -163 1463 -125
rect 1417 -197 1423 -163
rect 1457 -197 1463 -163
rect 1417 -235 1463 -197
rect 1417 -269 1423 -235
rect 1457 -269 1463 -235
rect 1417 -300 1463 -269
rect 1513 269 1559 300
rect 1513 235 1519 269
rect 1553 235 1559 269
rect 1513 197 1559 235
rect 1513 163 1519 197
rect 1553 163 1559 197
rect 1513 125 1559 163
rect 1513 91 1519 125
rect 1553 91 1559 125
rect 1513 53 1559 91
rect 1513 19 1519 53
rect 1553 19 1559 53
rect 1513 -19 1559 19
rect 1513 -53 1519 -19
rect 1553 -53 1559 -19
rect 1513 -91 1559 -53
rect 1513 -125 1519 -91
rect 1553 -125 1559 -91
rect 1513 -163 1559 -125
rect 1513 -197 1519 -163
rect 1553 -197 1559 -163
rect 1513 -235 1559 -197
rect 1513 -269 1519 -235
rect 1553 -269 1559 -235
rect 1513 -300 1559 -269
rect 1609 269 1655 300
rect 1609 235 1615 269
rect 1649 235 1655 269
rect 1609 197 1655 235
rect 1609 163 1615 197
rect 1649 163 1655 197
rect 1609 125 1655 163
rect 1609 91 1615 125
rect 1649 91 1655 125
rect 1609 53 1655 91
rect 1609 19 1615 53
rect 1649 19 1655 53
rect 1609 -19 1655 19
rect 1609 -53 1615 -19
rect 1649 -53 1655 -19
rect 1609 -91 1655 -53
rect 1609 -125 1615 -91
rect 1649 -125 1655 -91
rect 1609 -163 1655 -125
rect 1609 -197 1615 -163
rect 1649 -197 1655 -163
rect 1609 -235 1655 -197
rect 1609 -269 1615 -235
rect 1649 -269 1655 -235
rect 1609 -300 1655 -269
rect 1705 269 1751 300
rect 1705 235 1711 269
rect 1745 235 1751 269
rect 1705 197 1751 235
rect 1705 163 1711 197
rect 1745 163 1751 197
rect 1705 125 1751 163
rect 1705 91 1711 125
rect 1745 91 1751 125
rect 1705 53 1751 91
rect 1705 19 1711 53
rect 1745 19 1751 53
rect 1705 -19 1751 19
rect 1705 -53 1711 -19
rect 1745 -53 1751 -19
rect 1705 -91 1751 -53
rect 1705 -125 1711 -91
rect 1745 -125 1751 -91
rect 1705 -163 1751 -125
rect 1705 -197 1711 -163
rect 1745 -197 1751 -163
rect 1705 -235 1751 -197
rect 1705 -269 1711 -235
rect 1745 -269 1751 -235
rect 1705 -300 1751 -269
rect 1801 269 1847 300
rect 1801 235 1807 269
rect 1841 235 1847 269
rect 1801 197 1847 235
rect 1801 163 1807 197
rect 1841 163 1847 197
rect 1801 125 1847 163
rect 1801 91 1807 125
rect 1841 91 1847 125
rect 1801 53 1847 91
rect 1801 19 1807 53
rect 1841 19 1847 53
rect 1801 -19 1847 19
rect 1801 -53 1807 -19
rect 1841 -53 1847 -19
rect 1801 -91 1847 -53
rect 1801 -125 1807 -91
rect 1841 -125 1847 -91
rect 1801 -163 1847 -125
rect 1801 -197 1807 -163
rect 1841 -197 1847 -163
rect 1801 -235 1847 -197
rect 1801 -269 1807 -235
rect 1841 -269 1847 -235
rect 1801 -300 1847 -269
rect 1897 269 1943 300
rect 1897 235 1903 269
rect 1937 235 1943 269
rect 1897 197 1943 235
rect 1897 163 1903 197
rect 1937 163 1943 197
rect 1897 125 1943 163
rect 1897 91 1903 125
rect 1937 91 1943 125
rect 1897 53 1943 91
rect 1897 19 1903 53
rect 1937 19 1943 53
rect 1897 -19 1943 19
rect 1897 -53 1903 -19
rect 1937 -53 1943 -19
rect 1897 -91 1943 -53
rect 1897 -125 1903 -91
rect 1937 -125 1943 -91
rect 1897 -163 1943 -125
rect 1897 -197 1903 -163
rect 1937 -197 1943 -163
rect 1897 -235 1943 -197
rect 1897 -269 1903 -235
rect 1937 -269 1943 -235
rect 1897 -300 1943 -269
rect 1993 269 2039 300
rect 1993 235 1999 269
rect 2033 235 2039 269
rect 1993 197 2039 235
rect 1993 163 1999 197
rect 2033 163 2039 197
rect 1993 125 2039 163
rect 1993 91 1999 125
rect 2033 91 2039 125
rect 1993 53 2039 91
rect 1993 19 1999 53
rect 2033 19 2039 53
rect 1993 -19 2039 19
rect 1993 -53 1999 -19
rect 2033 -53 2039 -19
rect 1993 -91 2039 -53
rect 1993 -125 1999 -91
rect 2033 -125 2039 -91
rect 1993 -163 2039 -125
rect 1993 -197 1999 -163
rect 2033 -197 2039 -163
rect 1993 -235 2039 -197
rect 1993 -269 1999 -235
rect 2033 -269 2039 -235
rect 1993 -300 2039 -269
rect -1997 -338 -1939 -332
rect -1997 -372 -1985 -338
rect -1951 -372 -1939 -338
rect -1997 -378 -1939 -372
rect -1805 -338 -1747 -332
rect -1805 -372 -1793 -338
rect -1759 -372 -1747 -338
rect -1805 -378 -1747 -372
rect -1613 -338 -1555 -332
rect -1613 -372 -1601 -338
rect -1567 -372 -1555 -338
rect -1613 -378 -1555 -372
rect -1421 -338 -1363 -332
rect -1421 -372 -1409 -338
rect -1375 -372 -1363 -338
rect -1421 -378 -1363 -372
rect -1229 -338 -1171 -332
rect -1229 -372 -1217 -338
rect -1183 -372 -1171 -338
rect -1229 -378 -1171 -372
rect -1037 -338 -979 -332
rect -1037 -372 -1025 -338
rect -991 -372 -979 -338
rect -1037 -378 -979 -372
rect -845 -338 -787 -332
rect -845 -372 -833 -338
rect -799 -372 -787 -338
rect -845 -378 -787 -372
rect -653 -338 -595 -332
rect -653 -372 -641 -338
rect -607 -372 -595 -338
rect -653 -378 -595 -372
rect -461 -338 -403 -332
rect -461 -372 -449 -338
rect -415 -372 -403 -338
rect -461 -378 -403 -372
rect -269 -338 -211 -332
rect -269 -372 -257 -338
rect -223 -372 -211 -338
rect -269 -378 -211 -372
rect -77 -338 -19 -332
rect -77 -372 -65 -338
rect -31 -372 -19 -338
rect -77 -378 -19 -372
rect 115 -338 173 -332
rect 115 -372 127 -338
rect 161 -372 173 -338
rect 115 -378 173 -372
rect 307 -338 365 -332
rect 307 -372 319 -338
rect 353 -372 365 -338
rect 307 -378 365 -372
rect 499 -338 557 -332
rect 499 -372 511 -338
rect 545 -372 557 -338
rect 499 -378 557 -372
rect 691 -338 749 -332
rect 691 -372 703 -338
rect 737 -372 749 -338
rect 691 -378 749 -372
rect 883 -338 941 -332
rect 883 -372 895 -338
rect 929 -372 941 -338
rect 883 -378 941 -372
rect 1075 -338 1133 -332
rect 1075 -372 1087 -338
rect 1121 -372 1133 -338
rect 1075 -378 1133 -372
rect 1267 -338 1325 -332
rect 1267 -372 1279 -338
rect 1313 -372 1325 -338
rect 1267 -378 1325 -372
rect 1459 -338 1517 -332
rect 1459 -372 1471 -338
rect 1505 -372 1517 -338
rect 1459 -378 1517 -372
rect 1651 -338 1709 -332
rect 1651 -372 1663 -338
rect 1697 -372 1709 -338
rect 1651 -378 1709 -372
rect 1843 -338 1901 -332
rect 1843 -372 1855 -338
rect 1889 -372 1901 -338
rect 1843 -378 1901 -372
<< properties >>
string FIXED_BBOX -2130 -457 2130 457
<< end >>
