magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 535 35 967
rect -35 -967 35 -535
<< ppolyres >>
rect -35 -535 35 535
<< viali >>
rect -17 913 17 947
rect -17 841 17 875
rect -17 769 17 803
rect -17 697 17 731
rect -17 625 17 659
rect -17 553 17 587
rect -17 -588 17 -554
rect -17 -660 17 -626
rect -17 -732 17 -698
rect -17 -804 17 -770
rect -17 -876 17 -842
rect -17 -948 17 -914
<< metal1 >>
rect -25 947 25 961
rect -25 913 -17 947
rect 17 913 25 947
rect -25 875 25 913
rect -25 841 -17 875
rect 17 841 25 875
rect -25 803 25 841
rect -25 769 -17 803
rect 17 769 25 803
rect -25 731 25 769
rect -25 697 -17 731
rect 17 697 25 731
rect -25 659 25 697
rect -25 625 -17 659
rect 17 625 25 659
rect -25 587 25 625
rect -25 553 -17 587
rect 17 553 25 587
rect -25 540 25 553
rect -25 -554 25 -540
rect -25 -588 -17 -554
rect 17 -588 25 -554
rect -25 -626 25 -588
rect -25 -660 -17 -626
rect 17 -660 25 -626
rect -25 -698 25 -660
rect -25 -732 -17 -698
rect 17 -732 25 -698
rect -25 -770 25 -732
rect -25 -804 -17 -770
rect 17 -804 25 -770
rect -25 -842 25 -804
rect -25 -876 -17 -842
rect 17 -876 25 -842
rect -25 -914 25 -876
rect -25 -948 -17 -914
rect 17 -948 25 -914
rect -25 -961 25 -948
<< end >>
