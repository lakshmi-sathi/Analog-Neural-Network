magic
tech sky130A
magscale 1 2
timestamp 1626782926
<< error_p >>
rect -173 581 -115 587
rect 19 581 77 587
rect 211 581 269 587
rect -173 547 -161 581
rect 19 547 31 581
rect 211 547 223 581
rect -173 541 -115 547
rect 19 541 77 547
rect 211 541 269 547
rect -269 -547 -211 -541
rect -77 -547 -19 -541
rect 115 -547 173 -541
rect -269 -581 -257 -547
rect -77 -581 -65 -547
rect 115 -581 127 -547
rect -269 -587 -211 -581
rect -77 -587 -19 -581
rect 115 -587 173 -581
<< nwell >>
rect -455 -719 455 719
<< pmos >>
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
<< pdiff >>
rect -317 488 -255 500
rect -317 -488 -305 488
rect -271 -488 -255 488
rect -317 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 317 500
rect 255 -488 271 488
rect 305 -488 317 488
rect 255 -500 317 -488
<< pdiffc >>
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
<< nsubdiff >>
rect -419 649 -323 683
rect 323 649 419 683
rect -419 587 -385 649
rect 385 587 419 649
rect -419 -649 -385 -587
rect 385 -649 419 -587
rect -419 -683 -323 -649
rect 323 -683 419 -649
<< nsubdiffcont >>
rect -323 649 323 683
rect -419 -587 -385 587
rect 385 -587 419 587
rect -323 -683 323 -649
<< poly >>
rect -177 581 -111 597
rect -177 547 -161 581
rect -127 547 -111 581
rect -177 531 -111 547
rect 15 581 81 597
rect 15 547 31 581
rect 65 547 81 581
rect 15 531 81 547
rect 207 581 273 597
rect 207 547 223 581
rect 257 547 273 581
rect 207 531 273 547
rect -255 500 -225 526
rect -159 500 -129 531
rect -63 500 -33 526
rect 33 500 63 531
rect 129 500 159 526
rect 225 500 255 531
rect -255 -531 -225 -500
rect -159 -526 -129 -500
rect -63 -531 -33 -500
rect 33 -526 63 -500
rect 129 -531 159 -500
rect 225 -526 255 -500
rect -273 -547 -207 -531
rect -273 -581 -257 -547
rect -223 -581 -207 -547
rect -273 -597 -207 -581
rect -81 -547 -15 -531
rect -81 -581 -65 -547
rect -31 -581 -15 -547
rect -81 -597 -15 -581
rect 111 -547 177 -531
rect 111 -581 127 -547
rect 161 -581 177 -547
rect 111 -597 177 -581
<< polycont >>
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect -257 -581 -223 -547
rect -65 -581 -31 -547
rect 127 -581 161 -547
<< locali >>
rect -419 649 -323 683
rect 323 649 419 683
rect -419 587 -385 649
rect 385 587 419 649
rect -177 547 -161 581
rect -127 547 -111 581
rect 15 547 31 581
rect 65 547 81 581
rect 207 547 223 581
rect 257 547 273 581
rect -305 488 -271 504
rect -305 -504 -271 -488
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
rect 271 488 305 504
rect 271 -504 305 -488
rect -273 -581 -257 -547
rect -223 -581 -207 -547
rect -81 -581 -65 -547
rect -31 -581 -15 -547
rect 111 -581 127 -547
rect 161 -581 177 -547
rect -419 -649 -385 -587
rect 385 -649 419 -587
rect -419 -683 -323 -649
rect 323 -683 419 -649
<< viali >>
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect -257 -581 -223 -547
rect -65 -581 -31 -547
rect 127 -581 161 -547
<< metal1 >>
rect -173 581 -115 587
rect -173 547 -161 581
rect -127 547 -115 581
rect -173 541 -115 547
rect 19 581 77 587
rect 19 547 31 581
rect 65 547 77 581
rect 19 541 77 547
rect 211 581 269 587
rect 211 547 223 581
rect 257 547 269 581
rect 211 541 269 547
rect -311 488 -265 500
rect -311 -488 -305 488
rect -271 -488 -265 488
rect -311 -500 -265 -488
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect 265 488 311 500
rect 265 -488 271 488
rect 305 -488 311 488
rect 265 -500 311 -488
rect -269 -547 -211 -541
rect -269 -581 -257 -547
rect -223 -581 -211 -547
rect -269 -587 -211 -581
rect -77 -547 -19 -541
rect -77 -581 -65 -547
rect -31 -581 -19 -547
rect -77 -587 -19 -581
rect 115 -547 173 -541
rect 115 -581 127 -547
rect 161 -581 173 -547
rect 115 -587 173 -581
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -402 -666 402 666
string parameters w 5 l 0.15 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
