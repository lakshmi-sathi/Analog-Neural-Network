magic
tech sky130A
magscale 1 2
timestamp 1626793425
<< error_p >>
rect -269 1997 -211 2003
rect -77 1997 -19 2003
rect 115 1997 173 2003
rect -269 1963 -257 1997
rect -77 1963 -65 1997
rect 115 1963 127 1997
rect -269 1957 -211 1963
rect -77 1957 -19 1963
rect 115 1957 173 1963
rect -173 1427 -115 1433
rect 19 1427 77 1433
rect 211 1427 269 1433
rect -173 1393 -161 1427
rect 19 1393 31 1427
rect 211 1393 223 1427
rect -173 1387 -115 1393
rect 19 1387 77 1393
rect 211 1387 269 1393
rect -173 1319 -115 1325
rect 19 1319 77 1325
rect 211 1319 269 1325
rect -173 1285 -161 1319
rect 19 1285 31 1319
rect 211 1285 223 1319
rect -173 1279 -115 1285
rect 19 1279 77 1285
rect 211 1279 269 1285
rect -269 749 -211 755
rect -77 749 -19 755
rect 115 749 173 755
rect -269 715 -257 749
rect -77 715 -65 749
rect 115 715 127 749
rect -269 709 -211 715
rect -77 709 -19 715
rect 115 709 173 715
rect -269 641 -211 647
rect -77 641 -19 647
rect 115 641 173 647
rect -269 607 -257 641
rect -77 607 -65 641
rect 115 607 127 641
rect -269 601 -211 607
rect -77 601 -19 607
rect 115 601 173 607
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect -269 -607 -211 -601
rect -77 -607 -19 -601
rect 115 -607 173 -601
rect -269 -641 -257 -607
rect -77 -641 -65 -607
rect 115 -641 127 -607
rect -269 -647 -211 -641
rect -77 -647 -19 -641
rect 115 -647 173 -641
rect -269 -715 -211 -709
rect -77 -715 -19 -709
rect 115 -715 173 -709
rect -269 -749 -257 -715
rect -77 -749 -65 -715
rect 115 -749 127 -715
rect -269 -755 -211 -749
rect -77 -755 -19 -749
rect 115 -755 173 -749
rect -173 -1285 -115 -1279
rect 19 -1285 77 -1279
rect 211 -1285 269 -1279
rect -173 -1319 -161 -1285
rect 19 -1319 31 -1285
rect 211 -1319 223 -1285
rect -173 -1325 -115 -1319
rect 19 -1325 77 -1319
rect 211 -1325 269 -1319
rect -173 -1393 -115 -1387
rect 19 -1393 77 -1387
rect 211 -1393 269 -1387
rect -173 -1427 -161 -1393
rect 19 -1427 31 -1393
rect 211 -1427 223 -1393
rect -173 -1433 -115 -1427
rect 19 -1433 77 -1427
rect 211 -1433 269 -1427
rect -269 -1963 -211 -1957
rect -77 -1963 -19 -1957
rect 115 -1963 173 -1957
rect -269 -1997 -257 -1963
rect -77 -1997 -65 -1963
rect 115 -1997 127 -1963
rect -269 -2003 -211 -1997
rect -77 -2003 -19 -1997
rect 115 -2003 173 -1997
<< nwell >>
rect -455 -2135 455 2135
<< pmos >>
rect -255 1474 -225 1916
rect -159 1474 -129 1916
rect -63 1474 -33 1916
rect 33 1474 63 1916
rect 129 1474 159 1916
rect 225 1474 255 1916
rect -255 796 -225 1238
rect -159 796 -129 1238
rect -63 796 -33 1238
rect 33 796 63 1238
rect 129 796 159 1238
rect 225 796 255 1238
rect -255 118 -225 560
rect -159 118 -129 560
rect -63 118 -33 560
rect 33 118 63 560
rect 129 118 159 560
rect 225 118 255 560
rect -255 -560 -225 -118
rect -159 -560 -129 -118
rect -63 -560 -33 -118
rect 33 -560 63 -118
rect 129 -560 159 -118
rect 225 -560 255 -118
rect -255 -1238 -225 -796
rect -159 -1238 -129 -796
rect -63 -1238 -33 -796
rect 33 -1238 63 -796
rect 129 -1238 159 -796
rect 225 -1238 255 -796
rect -255 -1916 -225 -1474
rect -159 -1916 -129 -1474
rect -63 -1916 -33 -1474
rect 33 -1916 63 -1474
rect 129 -1916 159 -1474
rect 225 -1916 255 -1474
<< pdiff >>
rect -317 1904 -255 1916
rect -317 1486 -305 1904
rect -271 1486 -255 1904
rect -317 1474 -255 1486
rect -225 1904 -159 1916
rect -225 1486 -209 1904
rect -175 1486 -159 1904
rect -225 1474 -159 1486
rect -129 1904 -63 1916
rect -129 1486 -113 1904
rect -79 1486 -63 1904
rect -129 1474 -63 1486
rect -33 1904 33 1916
rect -33 1486 -17 1904
rect 17 1486 33 1904
rect -33 1474 33 1486
rect 63 1904 129 1916
rect 63 1486 79 1904
rect 113 1486 129 1904
rect 63 1474 129 1486
rect 159 1904 225 1916
rect 159 1486 175 1904
rect 209 1486 225 1904
rect 159 1474 225 1486
rect 255 1904 317 1916
rect 255 1486 271 1904
rect 305 1486 317 1904
rect 255 1474 317 1486
rect -317 1226 -255 1238
rect -317 808 -305 1226
rect -271 808 -255 1226
rect -317 796 -255 808
rect -225 1226 -159 1238
rect -225 808 -209 1226
rect -175 808 -159 1226
rect -225 796 -159 808
rect -129 1226 -63 1238
rect -129 808 -113 1226
rect -79 808 -63 1226
rect -129 796 -63 808
rect -33 1226 33 1238
rect -33 808 -17 1226
rect 17 808 33 1226
rect -33 796 33 808
rect 63 1226 129 1238
rect 63 808 79 1226
rect 113 808 129 1226
rect 63 796 129 808
rect 159 1226 225 1238
rect 159 808 175 1226
rect 209 808 225 1226
rect 159 796 225 808
rect 255 1226 317 1238
rect 255 808 271 1226
rect 305 808 317 1226
rect 255 796 317 808
rect -317 548 -255 560
rect -317 130 -305 548
rect -271 130 -255 548
rect -317 118 -255 130
rect -225 548 -159 560
rect -225 130 -209 548
rect -175 130 -159 548
rect -225 118 -159 130
rect -129 548 -63 560
rect -129 130 -113 548
rect -79 130 -63 548
rect -129 118 -63 130
rect -33 548 33 560
rect -33 130 -17 548
rect 17 130 33 548
rect -33 118 33 130
rect 63 548 129 560
rect 63 130 79 548
rect 113 130 129 548
rect 63 118 129 130
rect 159 548 225 560
rect 159 130 175 548
rect 209 130 225 548
rect 159 118 225 130
rect 255 548 317 560
rect 255 130 271 548
rect 305 130 317 548
rect 255 118 317 130
rect -317 -130 -255 -118
rect -317 -548 -305 -130
rect -271 -548 -255 -130
rect -317 -560 -255 -548
rect -225 -130 -159 -118
rect -225 -548 -209 -130
rect -175 -548 -159 -130
rect -225 -560 -159 -548
rect -129 -130 -63 -118
rect -129 -548 -113 -130
rect -79 -548 -63 -130
rect -129 -560 -63 -548
rect -33 -130 33 -118
rect -33 -548 -17 -130
rect 17 -548 33 -130
rect -33 -560 33 -548
rect 63 -130 129 -118
rect 63 -548 79 -130
rect 113 -548 129 -130
rect 63 -560 129 -548
rect 159 -130 225 -118
rect 159 -548 175 -130
rect 209 -548 225 -130
rect 159 -560 225 -548
rect 255 -130 317 -118
rect 255 -548 271 -130
rect 305 -548 317 -130
rect 255 -560 317 -548
rect -317 -808 -255 -796
rect -317 -1226 -305 -808
rect -271 -1226 -255 -808
rect -317 -1238 -255 -1226
rect -225 -808 -159 -796
rect -225 -1226 -209 -808
rect -175 -1226 -159 -808
rect -225 -1238 -159 -1226
rect -129 -808 -63 -796
rect -129 -1226 -113 -808
rect -79 -1226 -63 -808
rect -129 -1238 -63 -1226
rect -33 -808 33 -796
rect -33 -1226 -17 -808
rect 17 -1226 33 -808
rect -33 -1238 33 -1226
rect 63 -808 129 -796
rect 63 -1226 79 -808
rect 113 -1226 129 -808
rect 63 -1238 129 -1226
rect 159 -808 225 -796
rect 159 -1226 175 -808
rect 209 -1226 225 -808
rect 159 -1238 225 -1226
rect 255 -808 317 -796
rect 255 -1226 271 -808
rect 305 -1226 317 -808
rect 255 -1238 317 -1226
rect -317 -1486 -255 -1474
rect -317 -1904 -305 -1486
rect -271 -1904 -255 -1486
rect -317 -1916 -255 -1904
rect -225 -1486 -159 -1474
rect -225 -1904 -209 -1486
rect -175 -1904 -159 -1486
rect -225 -1916 -159 -1904
rect -129 -1486 -63 -1474
rect -129 -1904 -113 -1486
rect -79 -1904 -63 -1486
rect -129 -1916 -63 -1904
rect -33 -1486 33 -1474
rect -33 -1904 -17 -1486
rect 17 -1904 33 -1486
rect -33 -1916 33 -1904
rect 63 -1486 129 -1474
rect 63 -1904 79 -1486
rect 113 -1904 129 -1486
rect 63 -1916 129 -1904
rect 159 -1486 225 -1474
rect 159 -1904 175 -1486
rect 209 -1904 225 -1486
rect 159 -1916 225 -1904
rect 255 -1486 317 -1474
rect 255 -1904 271 -1486
rect 305 -1904 317 -1486
rect 255 -1916 317 -1904
<< pdiffc >>
rect -305 1486 -271 1904
rect -209 1486 -175 1904
rect -113 1486 -79 1904
rect -17 1486 17 1904
rect 79 1486 113 1904
rect 175 1486 209 1904
rect 271 1486 305 1904
rect -305 808 -271 1226
rect -209 808 -175 1226
rect -113 808 -79 1226
rect -17 808 17 1226
rect 79 808 113 1226
rect 175 808 209 1226
rect 271 808 305 1226
rect -305 130 -271 548
rect -209 130 -175 548
rect -113 130 -79 548
rect -17 130 17 548
rect 79 130 113 548
rect 175 130 209 548
rect 271 130 305 548
rect -305 -548 -271 -130
rect -209 -548 -175 -130
rect -113 -548 -79 -130
rect -17 -548 17 -130
rect 79 -548 113 -130
rect 175 -548 209 -130
rect 271 -548 305 -130
rect -305 -1226 -271 -808
rect -209 -1226 -175 -808
rect -113 -1226 -79 -808
rect -17 -1226 17 -808
rect 79 -1226 113 -808
rect 175 -1226 209 -808
rect 271 -1226 305 -808
rect -305 -1904 -271 -1486
rect -209 -1904 -175 -1486
rect -113 -1904 -79 -1486
rect -17 -1904 17 -1486
rect 79 -1904 113 -1486
rect 175 -1904 209 -1486
rect 271 -1904 305 -1486
<< nsubdiff >>
rect -419 2065 -323 2099
rect 323 2065 419 2099
rect -419 2003 -385 2065
rect 385 2003 419 2065
rect -419 -2065 -385 -2003
rect 385 -2065 419 -2003
rect -419 -2099 -323 -2065
rect 323 -2099 419 -2065
<< nsubdiffcont >>
rect -323 2065 323 2099
rect -419 -2003 -385 2003
rect 385 -2003 419 2003
rect -323 -2099 323 -2065
<< poly >>
rect -273 1997 -207 2013
rect -273 1963 -257 1997
rect -223 1963 -207 1997
rect -273 1947 -207 1963
rect -81 1997 -15 2013
rect -81 1963 -65 1997
rect -31 1963 -15 1997
rect -81 1947 -15 1963
rect 111 1997 177 2013
rect 111 1963 127 1997
rect 161 1963 177 1997
rect 111 1947 177 1963
rect -255 1916 -225 1947
rect -159 1916 -129 1942
rect -63 1916 -33 1947
rect 33 1916 63 1942
rect 129 1916 159 1947
rect 225 1916 255 1942
rect -255 1448 -225 1474
rect -159 1443 -129 1474
rect -63 1448 -33 1474
rect 33 1443 63 1474
rect 129 1448 159 1474
rect 225 1443 255 1474
rect -177 1427 -111 1443
rect -177 1393 -161 1427
rect -127 1393 -111 1427
rect -177 1377 -111 1393
rect 15 1427 81 1443
rect 15 1393 31 1427
rect 65 1393 81 1427
rect 15 1377 81 1393
rect 207 1427 273 1443
rect 207 1393 223 1427
rect 257 1393 273 1427
rect 207 1377 273 1393
rect -177 1319 -111 1335
rect -177 1285 -161 1319
rect -127 1285 -111 1319
rect -177 1269 -111 1285
rect 15 1319 81 1335
rect 15 1285 31 1319
rect 65 1285 81 1319
rect 15 1269 81 1285
rect 207 1319 273 1335
rect 207 1285 223 1319
rect 257 1285 273 1319
rect 207 1269 273 1285
rect -255 1238 -225 1264
rect -159 1238 -129 1269
rect -63 1238 -33 1264
rect 33 1238 63 1269
rect 129 1238 159 1264
rect 225 1238 255 1269
rect -255 765 -225 796
rect -159 770 -129 796
rect -63 765 -33 796
rect 33 770 63 796
rect 129 765 159 796
rect 225 770 255 796
rect -273 749 -207 765
rect -273 715 -257 749
rect -223 715 -207 749
rect -273 699 -207 715
rect -81 749 -15 765
rect -81 715 -65 749
rect -31 715 -15 749
rect -81 699 -15 715
rect 111 749 177 765
rect 111 715 127 749
rect 161 715 177 749
rect 111 699 177 715
rect -273 641 -207 657
rect -273 607 -257 641
rect -223 607 -207 641
rect -273 591 -207 607
rect -81 641 -15 657
rect -81 607 -65 641
rect -31 607 -15 641
rect -81 591 -15 607
rect 111 641 177 657
rect 111 607 127 641
rect 161 607 177 641
rect 111 591 177 607
rect -255 560 -225 591
rect -159 560 -129 586
rect -63 560 -33 591
rect 33 560 63 586
rect 129 560 159 591
rect 225 560 255 586
rect -255 92 -225 118
rect -159 87 -129 118
rect -63 92 -33 118
rect 33 87 63 118
rect 129 92 159 118
rect 225 87 255 118
rect -177 71 -111 87
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 207 -87 273 -71
rect -255 -118 -225 -92
rect -159 -118 -129 -87
rect -63 -118 -33 -92
rect 33 -118 63 -87
rect 129 -118 159 -92
rect 225 -118 255 -87
rect -255 -591 -225 -560
rect -159 -586 -129 -560
rect -63 -591 -33 -560
rect 33 -586 63 -560
rect 129 -591 159 -560
rect 225 -586 255 -560
rect -273 -607 -207 -591
rect -273 -641 -257 -607
rect -223 -641 -207 -607
rect -273 -657 -207 -641
rect -81 -607 -15 -591
rect -81 -641 -65 -607
rect -31 -641 -15 -607
rect -81 -657 -15 -641
rect 111 -607 177 -591
rect 111 -641 127 -607
rect 161 -641 177 -607
rect 111 -657 177 -641
rect -273 -715 -207 -699
rect -273 -749 -257 -715
rect -223 -749 -207 -715
rect -273 -765 -207 -749
rect -81 -715 -15 -699
rect -81 -749 -65 -715
rect -31 -749 -15 -715
rect -81 -765 -15 -749
rect 111 -715 177 -699
rect 111 -749 127 -715
rect 161 -749 177 -715
rect 111 -765 177 -749
rect -255 -796 -225 -765
rect -159 -796 -129 -770
rect -63 -796 -33 -765
rect 33 -796 63 -770
rect 129 -796 159 -765
rect 225 -796 255 -770
rect -255 -1264 -225 -1238
rect -159 -1269 -129 -1238
rect -63 -1264 -33 -1238
rect 33 -1269 63 -1238
rect 129 -1264 159 -1238
rect 225 -1269 255 -1238
rect -177 -1285 -111 -1269
rect -177 -1319 -161 -1285
rect -127 -1319 -111 -1285
rect -177 -1335 -111 -1319
rect 15 -1285 81 -1269
rect 15 -1319 31 -1285
rect 65 -1319 81 -1285
rect 15 -1335 81 -1319
rect 207 -1285 273 -1269
rect 207 -1319 223 -1285
rect 257 -1319 273 -1285
rect 207 -1335 273 -1319
rect -177 -1393 -111 -1377
rect -177 -1427 -161 -1393
rect -127 -1427 -111 -1393
rect -177 -1443 -111 -1427
rect 15 -1393 81 -1377
rect 15 -1427 31 -1393
rect 65 -1427 81 -1393
rect 15 -1443 81 -1427
rect 207 -1393 273 -1377
rect 207 -1427 223 -1393
rect 257 -1427 273 -1393
rect 207 -1443 273 -1427
rect -255 -1474 -225 -1448
rect -159 -1474 -129 -1443
rect -63 -1474 -33 -1448
rect 33 -1474 63 -1443
rect 129 -1474 159 -1448
rect 225 -1474 255 -1443
rect -255 -1947 -225 -1916
rect -159 -1942 -129 -1916
rect -63 -1947 -33 -1916
rect 33 -1942 63 -1916
rect 129 -1947 159 -1916
rect 225 -1942 255 -1916
rect -273 -1963 -207 -1947
rect -273 -1997 -257 -1963
rect -223 -1997 -207 -1963
rect -273 -2013 -207 -1997
rect -81 -1963 -15 -1947
rect -81 -1997 -65 -1963
rect -31 -1997 -15 -1963
rect -81 -2013 -15 -1997
rect 111 -1963 177 -1947
rect 111 -1997 127 -1963
rect 161 -1997 177 -1963
rect 111 -2013 177 -1997
<< polycont >>
rect -257 1963 -223 1997
rect -65 1963 -31 1997
rect 127 1963 161 1997
rect -161 1393 -127 1427
rect 31 1393 65 1427
rect 223 1393 257 1427
rect -161 1285 -127 1319
rect 31 1285 65 1319
rect 223 1285 257 1319
rect -257 715 -223 749
rect -65 715 -31 749
rect 127 715 161 749
rect -257 607 -223 641
rect -65 607 -31 641
rect 127 607 161 641
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect -257 -641 -223 -607
rect -65 -641 -31 -607
rect 127 -641 161 -607
rect -257 -749 -223 -715
rect -65 -749 -31 -715
rect 127 -749 161 -715
rect -161 -1319 -127 -1285
rect 31 -1319 65 -1285
rect 223 -1319 257 -1285
rect -161 -1427 -127 -1393
rect 31 -1427 65 -1393
rect 223 -1427 257 -1393
rect -257 -1997 -223 -1963
rect -65 -1997 -31 -1963
rect 127 -1997 161 -1963
<< locali >>
rect -419 2065 -323 2099
rect 323 2065 419 2099
rect -419 2003 -385 2065
rect 385 2003 419 2065
rect -273 1963 -257 1997
rect -223 1963 -207 1997
rect -81 1963 -65 1997
rect -31 1963 -15 1997
rect 111 1963 127 1997
rect 161 1963 177 1997
rect -305 1904 -271 1920
rect -305 1470 -271 1486
rect -209 1904 -175 1920
rect -209 1470 -175 1486
rect -113 1904 -79 1920
rect -113 1470 -79 1486
rect -17 1904 17 1920
rect -17 1470 17 1486
rect 79 1904 113 1920
rect 79 1470 113 1486
rect 175 1904 209 1920
rect 175 1470 209 1486
rect 271 1904 305 1920
rect 271 1470 305 1486
rect -177 1393 -161 1427
rect -127 1393 -111 1427
rect 15 1393 31 1427
rect 65 1393 81 1427
rect 207 1393 223 1427
rect 257 1393 273 1427
rect -177 1285 -161 1319
rect -127 1285 -111 1319
rect 15 1285 31 1319
rect 65 1285 81 1319
rect 207 1285 223 1319
rect 257 1285 273 1319
rect -305 1226 -271 1242
rect -305 792 -271 808
rect -209 1226 -175 1242
rect -209 792 -175 808
rect -113 1226 -79 1242
rect -113 792 -79 808
rect -17 1226 17 1242
rect -17 792 17 808
rect 79 1226 113 1242
rect 79 792 113 808
rect 175 1226 209 1242
rect 175 792 209 808
rect 271 1226 305 1242
rect 271 792 305 808
rect -273 715 -257 749
rect -223 715 -207 749
rect -81 715 -65 749
rect -31 715 -15 749
rect 111 715 127 749
rect 161 715 177 749
rect -273 607 -257 641
rect -223 607 -207 641
rect -81 607 -65 641
rect -31 607 -15 641
rect 111 607 127 641
rect 161 607 177 641
rect -305 548 -271 564
rect -305 114 -271 130
rect -209 548 -175 564
rect -209 114 -175 130
rect -113 548 -79 564
rect -113 114 -79 130
rect -17 548 17 564
rect -17 114 17 130
rect 79 548 113 564
rect 79 114 113 130
rect 175 548 209 564
rect 175 114 209 130
rect 271 548 305 564
rect 271 114 305 130
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect -305 -130 -271 -114
rect -305 -564 -271 -548
rect -209 -130 -175 -114
rect -209 -564 -175 -548
rect -113 -130 -79 -114
rect -113 -564 -79 -548
rect -17 -130 17 -114
rect -17 -564 17 -548
rect 79 -130 113 -114
rect 79 -564 113 -548
rect 175 -130 209 -114
rect 175 -564 209 -548
rect 271 -130 305 -114
rect 271 -564 305 -548
rect -273 -641 -257 -607
rect -223 -641 -207 -607
rect -81 -641 -65 -607
rect -31 -641 -15 -607
rect 111 -641 127 -607
rect 161 -641 177 -607
rect -273 -749 -257 -715
rect -223 -749 -207 -715
rect -81 -749 -65 -715
rect -31 -749 -15 -715
rect 111 -749 127 -715
rect 161 -749 177 -715
rect -305 -808 -271 -792
rect -305 -1242 -271 -1226
rect -209 -808 -175 -792
rect -209 -1242 -175 -1226
rect -113 -808 -79 -792
rect -113 -1242 -79 -1226
rect -17 -808 17 -792
rect -17 -1242 17 -1226
rect 79 -808 113 -792
rect 79 -1242 113 -1226
rect 175 -808 209 -792
rect 175 -1242 209 -1226
rect 271 -808 305 -792
rect 271 -1242 305 -1226
rect -177 -1319 -161 -1285
rect -127 -1319 -111 -1285
rect 15 -1319 31 -1285
rect 65 -1319 81 -1285
rect 207 -1319 223 -1285
rect 257 -1319 273 -1285
rect -177 -1427 -161 -1393
rect -127 -1427 -111 -1393
rect 15 -1427 31 -1393
rect 65 -1427 81 -1393
rect 207 -1427 223 -1393
rect 257 -1427 273 -1393
rect -305 -1486 -271 -1470
rect -305 -1920 -271 -1904
rect -209 -1486 -175 -1470
rect -209 -1920 -175 -1904
rect -113 -1486 -79 -1470
rect -113 -1920 -79 -1904
rect -17 -1486 17 -1470
rect -17 -1920 17 -1904
rect 79 -1486 113 -1470
rect 79 -1920 113 -1904
rect 175 -1486 209 -1470
rect 175 -1920 209 -1904
rect 271 -1486 305 -1470
rect 271 -1920 305 -1904
rect -273 -1997 -257 -1963
rect -223 -1997 -207 -1963
rect -81 -1997 -65 -1963
rect -31 -1997 -15 -1963
rect 111 -1997 127 -1963
rect 161 -1997 177 -1963
rect -419 -2065 -385 -2003
rect 385 -2065 419 -2003
rect -419 -2099 -323 -2065
rect 323 -2099 419 -2065
<< viali >>
rect -257 1963 -223 1997
rect -65 1963 -31 1997
rect 127 1963 161 1997
rect -305 1486 -271 1904
rect -209 1486 -175 1904
rect -113 1486 -79 1904
rect -17 1486 17 1904
rect 79 1486 113 1904
rect 175 1486 209 1904
rect 271 1486 305 1904
rect -161 1393 -127 1427
rect 31 1393 65 1427
rect 223 1393 257 1427
rect -161 1285 -127 1319
rect 31 1285 65 1319
rect 223 1285 257 1319
rect -305 808 -271 1226
rect -209 808 -175 1226
rect -113 808 -79 1226
rect -17 808 17 1226
rect 79 808 113 1226
rect 175 808 209 1226
rect 271 808 305 1226
rect -257 715 -223 749
rect -65 715 -31 749
rect 127 715 161 749
rect -257 607 -223 641
rect -65 607 -31 641
rect 127 607 161 641
rect -305 130 -271 548
rect -209 130 -175 548
rect -113 130 -79 548
rect -17 130 17 548
rect 79 130 113 548
rect 175 130 209 548
rect 271 130 305 548
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect -305 -548 -271 -130
rect -209 -548 -175 -130
rect -113 -548 -79 -130
rect -17 -548 17 -130
rect 79 -548 113 -130
rect 175 -548 209 -130
rect 271 -548 305 -130
rect -257 -641 -223 -607
rect -65 -641 -31 -607
rect 127 -641 161 -607
rect -257 -749 -223 -715
rect -65 -749 -31 -715
rect 127 -749 161 -715
rect -305 -1226 -271 -808
rect -209 -1226 -175 -808
rect -113 -1226 -79 -808
rect -17 -1226 17 -808
rect 79 -1226 113 -808
rect 175 -1226 209 -808
rect 271 -1226 305 -808
rect -161 -1319 -127 -1285
rect 31 -1319 65 -1285
rect 223 -1319 257 -1285
rect -161 -1427 -127 -1393
rect 31 -1427 65 -1393
rect 223 -1427 257 -1393
rect -305 -1904 -271 -1486
rect -209 -1904 -175 -1486
rect -113 -1904 -79 -1486
rect -17 -1904 17 -1486
rect 79 -1904 113 -1486
rect 175 -1904 209 -1486
rect 271 -1904 305 -1486
rect -257 -1997 -223 -1963
rect -65 -1997 -31 -1963
rect 127 -1997 161 -1963
<< metal1 >>
rect -269 1997 -211 2003
rect -269 1963 -257 1997
rect -223 1963 -211 1997
rect -269 1957 -211 1963
rect -77 1997 -19 2003
rect -77 1963 -65 1997
rect -31 1963 -19 1997
rect -77 1957 -19 1963
rect 115 1997 173 2003
rect 115 1963 127 1997
rect 161 1963 173 1997
rect 115 1957 173 1963
rect -311 1904 -265 1916
rect -311 1486 -305 1904
rect -271 1486 -265 1904
rect -311 1474 -265 1486
rect -215 1904 -169 1916
rect -215 1486 -209 1904
rect -175 1486 -169 1904
rect -215 1474 -169 1486
rect -119 1904 -73 1916
rect -119 1486 -113 1904
rect -79 1486 -73 1904
rect -119 1474 -73 1486
rect -23 1904 23 1916
rect -23 1486 -17 1904
rect 17 1486 23 1904
rect -23 1474 23 1486
rect 73 1904 119 1916
rect 73 1486 79 1904
rect 113 1486 119 1904
rect 73 1474 119 1486
rect 169 1904 215 1916
rect 169 1486 175 1904
rect 209 1486 215 1904
rect 169 1474 215 1486
rect 265 1904 311 1916
rect 265 1486 271 1904
rect 305 1486 311 1904
rect 265 1474 311 1486
rect -173 1427 -115 1433
rect -173 1393 -161 1427
rect -127 1393 -115 1427
rect -173 1387 -115 1393
rect 19 1427 77 1433
rect 19 1393 31 1427
rect 65 1393 77 1427
rect 19 1387 77 1393
rect 211 1427 269 1433
rect 211 1393 223 1427
rect 257 1393 269 1427
rect 211 1387 269 1393
rect -173 1319 -115 1325
rect -173 1285 -161 1319
rect -127 1285 -115 1319
rect -173 1279 -115 1285
rect 19 1319 77 1325
rect 19 1285 31 1319
rect 65 1285 77 1319
rect 19 1279 77 1285
rect 211 1319 269 1325
rect 211 1285 223 1319
rect 257 1285 269 1319
rect 211 1279 269 1285
rect -311 1226 -265 1238
rect -311 808 -305 1226
rect -271 808 -265 1226
rect -311 796 -265 808
rect -215 1226 -169 1238
rect -215 808 -209 1226
rect -175 808 -169 1226
rect -215 796 -169 808
rect -119 1226 -73 1238
rect -119 808 -113 1226
rect -79 808 -73 1226
rect -119 796 -73 808
rect -23 1226 23 1238
rect -23 808 -17 1226
rect 17 808 23 1226
rect -23 796 23 808
rect 73 1226 119 1238
rect 73 808 79 1226
rect 113 808 119 1226
rect 73 796 119 808
rect 169 1226 215 1238
rect 169 808 175 1226
rect 209 808 215 1226
rect 169 796 215 808
rect 265 1226 311 1238
rect 265 808 271 1226
rect 305 808 311 1226
rect 265 796 311 808
rect -269 749 -211 755
rect -269 715 -257 749
rect -223 715 -211 749
rect -269 709 -211 715
rect -77 749 -19 755
rect -77 715 -65 749
rect -31 715 -19 749
rect -77 709 -19 715
rect 115 749 173 755
rect 115 715 127 749
rect 161 715 173 749
rect 115 709 173 715
rect -269 641 -211 647
rect -269 607 -257 641
rect -223 607 -211 641
rect -269 601 -211 607
rect -77 641 -19 647
rect -77 607 -65 641
rect -31 607 -19 641
rect -77 601 -19 607
rect 115 641 173 647
rect 115 607 127 641
rect 161 607 173 641
rect 115 601 173 607
rect -311 548 -265 560
rect -311 130 -305 548
rect -271 130 -265 548
rect -311 118 -265 130
rect -215 548 -169 560
rect -215 130 -209 548
rect -175 130 -169 548
rect -215 118 -169 130
rect -119 548 -73 560
rect -119 130 -113 548
rect -79 130 -73 548
rect -119 118 -73 130
rect -23 548 23 560
rect -23 130 -17 548
rect 17 130 23 548
rect -23 118 23 130
rect 73 548 119 560
rect 73 130 79 548
rect 113 130 119 548
rect 73 118 119 130
rect 169 548 215 560
rect 169 130 175 548
rect 209 130 215 548
rect 169 118 215 130
rect 265 548 311 560
rect 265 130 271 548
rect 305 130 311 548
rect 265 118 311 130
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect -311 -130 -265 -118
rect -311 -548 -305 -130
rect -271 -548 -265 -130
rect -311 -560 -265 -548
rect -215 -130 -169 -118
rect -215 -548 -209 -130
rect -175 -548 -169 -130
rect -215 -560 -169 -548
rect -119 -130 -73 -118
rect -119 -548 -113 -130
rect -79 -548 -73 -130
rect -119 -560 -73 -548
rect -23 -130 23 -118
rect -23 -548 -17 -130
rect 17 -548 23 -130
rect -23 -560 23 -548
rect 73 -130 119 -118
rect 73 -548 79 -130
rect 113 -548 119 -130
rect 73 -560 119 -548
rect 169 -130 215 -118
rect 169 -548 175 -130
rect 209 -548 215 -130
rect 169 -560 215 -548
rect 265 -130 311 -118
rect 265 -548 271 -130
rect 305 -548 311 -130
rect 265 -560 311 -548
rect -269 -607 -211 -601
rect -269 -641 -257 -607
rect -223 -641 -211 -607
rect -269 -647 -211 -641
rect -77 -607 -19 -601
rect -77 -641 -65 -607
rect -31 -641 -19 -607
rect -77 -647 -19 -641
rect 115 -607 173 -601
rect 115 -641 127 -607
rect 161 -641 173 -607
rect 115 -647 173 -641
rect -269 -715 -211 -709
rect -269 -749 -257 -715
rect -223 -749 -211 -715
rect -269 -755 -211 -749
rect -77 -715 -19 -709
rect -77 -749 -65 -715
rect -31 -749 -19 -715
rect -77 -755 -19 -749
rect 115 -715 173 -709
rect 115 -749 127 -715
rect 161 -749 173 -715
rect 115 -755 173 -749
rect -311 -808 -265 -796
rect -311 -1226 -305 -808
rect -271 -1226 -265 -808
rect -311 -1238 -265 -1226
rect -215 -808 -169 -796
rect -215 -1226 -209 -808
rect -175 -1226 -169 -808
rect -215 -1238 -169 -1226
rect -119 -808 -73 -796
rect -119 -1226 -113 -808
rect -79 -1226 -73 -808
rect -119 -1238 -73 -1226
rect -23 -808 23 -796
rect -23 -1226 -17 -808
rect 17 -1226 23 -808
rect -23 -1238 23 -1226
rect 73 -808 119 -796
rect 73 -1226 79 -808
rect 113 -1226 119 -808
rect 73 -1238 119 -1226
rect 169 -808 215 -796
rect 169 -1226 175 -808
rect 209 -1226 215 -808
rect 169 -1238 215 -1226
rect 265 -808 311 -796
rect 265 -1226 271 -808
rect 305 -1226 311 -808
rect 265 -1238 311 -1226
rect -173 -1285 -115 -1279
rect -173 -1319 -161 -1285
rect -127 -1319 -115 -1285
rect -173 -1325 -115 -1319
rect 19 -1285 77 -1279
rect 19 -1319 31 -1285
rect 65 -1319 77 -1285
rect 19 -1325 77 -1319
rect 211 -1285 269 -1279
rect 211 -1319 223 -1285
rect 257 -1319 269 -1285
rect 211 -1325 269 -1319
rect -173 -1393 -115 -1387
rect -173 -1427 -161 -1393
rect -127 -1427 -115 -1393
rect -173 -1433 -115 -1427
rect 19 -1393 77 -1387
rect 19 -1427 31 -1393
rect 65 -1427 77 -1393
rect 19 -1433 77 -1427
rect 211 -1393 269 -1387
rect 211 -1427 223 -1393
rect 257 -1427 269 -1393
rect 211 -1433 269 -1427
rect -311 -1486 -265 -1474
rect -311 -1904 -305 -1486
rect -271 -1904 -265 -1486
rect -311 -1916 -265 -1904
rect -215 -1486 -169 -1474
rect -215 -1904 -209 -1486
rect -175 -1904 -169 -1486
rect -215 -1916 -169 -1904
rect -119 -1486 -73 -1474
rect -119 -1904 -113 -1486
rect -79 -1904 -73 -1486
rect -119 -1916 -73 -1904
rect -23 -1486 23 -1474
rect -23 -1904 -17 -1486
rect 17 -1904 23 -1486
rect -23 -1916 23 -1904
rect 73 -1486 119 -1474
rect 73 -1904 79 -1486
rect 113 -1904 119 -1486
rect 73 -1916 119 -1904
rect 169 -1486 215 -1474
rect 169 -1904 175 -1486
rect 209 -1904 215 -1486
rect 169 -1916 215 -1904
rect 265 -1486 311 -1474
rect 265 -1904 271 -1486
rect 305 -1904 311 -1486
rect 265 -1916 311 -1904
rect -269 -1963 -211 -1957
rect -269 -1997 -257 -1963
rect -223 -1997 -211 -1963
rect -269 -2003 -211 -1997
rect -77 -1963 -19 -1957
rect -77 -1997 -65 -1963
rect -31 -1997 -19 -1963
rect -77 -2003 -19 -1997
rect 115 -1963 173 -1957
rect 115 -1997 127 -1963
rect 161 -1997 173 -1963
rect 115 -2003 173 -1997
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -402 -2082 402 2082
string parameters w 2.21 l 0.15 m 6 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
