magic
tech sky130A
magscale 1 2
timestamp 1628069291
<< error_p >>
rect -269 521 -211 527
rect -77 521 -19 527
rect 115 521 173 527
rect 307 521 365 527
rect -269 487 -257 521
rect -77 487 -65 521
rect 115 487 127 521
rect 307 487 319 521
rect -269 481 -211 487
rect -77 481 -19 487
rect 115 481 173 487
rect 307 481 365 487
rect -365 -487 -307 -481
rect -173 -487 -115 -481
rect 19 -487 77 -481
rect 211 -487 269 -481
rect -365 -521 -353 -487
rect -173 -521 -161 -487
rect 19 -521 31 -487
rect 211 -521 223 -487
rect -365 -527 -307 -521
rect -173 -527 -115 -521
rect 19 -527 77 -521
rect 211 -527 269 -521
<< nwell >>
rect -551 -659 551 659
<< pmos >>
rect -351 -440 -321 440
rect -255 -440 -225 440
rect -159 -440 -129 440
rect -63 -440 -33 440
rect 33 -440 63 440
rect 129 -440 159 440
rect 225 -440 255 440
rect 321 -440 351 440
<< pdiff >>
rect -413 428 -351 440
rect -413 -428 -401 428
rect -367 -428 -351 428
rect -413 -440 -351 -428
rect -321 428 -255 440
rect -321 -428 -305 428
rect -271 -428 -255 428
rect -321 -440 -255 -428
rect -225 428 -159 440
rect -225 -428 -209 428
rect -175 -428 -159 428
rect -225 -440 -159 -428
rect -129 428 -63 440
rect -129 -428 -113 428
rect -79 -428 -63 428
rect -129 -440 -63 -428
rect -33 428 33 440
rect -33 -428 -17 428
rect 17 -428 33 428
rect -33 -440 33 -428
rect 63 428 129 440
rect 63 -428 79 428
rect 113 -428 129 428
rect 63 -440 129 -428
rect 159 428 225 440
rect 159 -428 175 428
rect 209 -428 225 428
rect 159 -440 225 -428
rect 255 428 321 440
rect 255 -428 271 428
rect 305 -428 321 428
rect 255 -440 321 -428
rect 351 428 413 440
rect 351 -428 367 428
rect 401 -428 413 428
rect 351 -440 413 -428
<< pdiffc >>
rect -401 -428 -367 428
rect -305 -428 -271 428
rect -209 -428 -175 428
rect -113 -428 -79 428
rect -17 -428 17 428
rect 79 -428 113 428
rect 175 -428 209 428
rect 271 -428 305 428
rect 367 -428 401 428
<< nsubdiff >>
rect -515 589 -419 623
rect 419 589 515 623
rect -515 527 -481 589
rect 481 527 515 589
rect -515 -589 -481 -527
rect 481 -589 515 -527
rect -515 -623 -419 -589
rect 419 -623 515 -589
<< nsubdiffcont >>
rect -419 589 419 623
rect -515 -527 -481 527
rect 481 -527 515 527
rect -419 -623 419 -589
<< poly >>
rect -273 521 -207 537
rect -273 487 -257 521
rect -223 487 -207 521
rect -273 471 -207 487
rect -81 521 -15 537
rect -81 487 -65 521
rect -31 487 -15 521
rect -81 471 -15 487
rect 111 521 177 537
rect 111 487 127 521
rect 161 487 177 521
rect 111 471 177 487
rect 303 521 369 537
rect 303 487 319 521
rect 353 487 369 521
rect 303 471 369 487
rect -351 440 -321 466
rect -255 440 -225 471
rect -159 440 -129 466
rect -63 440 -33 471
rect 33 440 63 466
rect 129 440 159 471
rect 225 440 255 466
rect 321 440 351 471
rect -351 -471 -321 -440
rect -255 -466 -225 -440
rect -159 -471 -129 -440
rect -63 -466 -33 -440
rect 33 -471 63 -440
rect 129 -466 159 -440
rect 225 -471 255 -440
rect 321 -466 351 -440
rect -369 -487 -303 -471
rect -369 -521 -353 -487
rect -319 -521 -303 -487
rect -369 -537 -303 -521
rect -177 -487 -111 -471
rect -177 -521 -161 -487
rect -127 -521 -111 -487
rect -177 -537 -111 -521
rect 15 -487 81 -471
rect 15 -521 31 -487
rect 65 -521 81 -487
rect 15 -537 81 -521
rect 207 -487 273 -471
rect 207 -521 223 -487
rect 257 -521 273 -487
rect 207 -537 273 -521
<< polycont >>
rect -257 487 -223 521
rect -65 487 -31 521
rect 127 487 161 521
rect 319 487 353 521
rect -353 -521 -319 -487
rect -161 -521 -127 -487
rect 31 -521 65 -487
rect 223 -521 257 -487
<< locali >>
rect -515 589 -419 623
rect 419 589 515 623
rect -515 527 -481 589
rect 481 527 515 589
rect -273 487 -257 521
rect -223 487 -207 521
rect -81 487 -65 521
rect -31 487 -15 521
rect 111 487 127 521
rect 161 487 177 521
rect 303 487 319 521
rect 353 487 369 521
rect -401 428 -367 444
rect -401 -444 -367 -428
rect -305 428 -271 444
rect -305 -444 -271 -428
rect -209 428 -175 444
rect -209 -444 -175 -428
rect -113 428 -79 444
rect -113 -444 -79 -428
rect -17 428 17 444
rect -17 -444 17 -428
rect 79 428 113 444
rect 79 -444 113 -428
rect 175 428 209 444
rect 175 -444 209 -428
rect 271 428 305 444
rect 271 -444 305 -428
rect 367 428 401 444
rect 367 -444 401 -428
rect -369 -521 -353 -487
rect -319 -521 -303 -487
rect -177 -521 -161 -487
rect -127 -521 -111 -487
rect 15 -521 31 -487
rect 65 -521 81 -487
rect 207 -521 223 -487
rect 257 -521 273 -487
rect -515 -589 -481 -527
rect 481 -589 515 -527
rect -515 -623 -419 -589
rect 419 -623 515 -589
<< viali >>
rect -257 487 -223 521
rect -65 487 -31 521
rect 127 487 161 521
rect 319 487 353 521
rect -401 -428 -367 428
rect -305 -428 -271 428
rect -209 -428 -175 428
rect -113 -428 -79 428
rect -17 -428 17 428
rect 79 -428 113 428
rect 175 -428 209 428
rect 271 -428 305 428
rect 367 -428 401 428
rect -353 -521 -319 -487
rect -161 -521 -127 -487
rect 31 -521 65 -487
rect 223 -521 257 -487
<< metal1 >>
rect -269 521 -211 527
rect -269 487 -257 521
rect -223 487 -211 521
rect -269 481 -211 487
rect -77 521 -19 527
rect -77 487 -65 521
rect -31 487 -19 521
rect -77 481 -19 487
rect 115 521 173 527
rect 115 487 127 521
rect 161 487 173 521
rect 115 481 173 487
rect 307 521 365 527
rect 307 487 319 521
rect 353 487 365 521
rect 307 481 365 487
rect -407 428 -361 440
rect -407 -428 -401 428
rect -367 -428 -361 428
rect -407 -440 -361 -428
rect -311 428 -265 440
rect -311 -428 -305 428
rect -271 -428 -265 428
rect -311 -440 -265 -428
rect -215 428 -169 440
rect -215 -428 -209 428
rect -175 -428 -169 428
rect -215 -440 -169 -428
rect -119 428 -73 440
rect -119 -428 -113 428
rect -79 -428 -73 428
rect -119 -440 -73 -428
rect -23 428 23 440
rect -23 -428 -17 428
rect 17 -428 23 428
rect -23 -440 23 -428
rect 73 428 119 440
rect 73 -428 79 428
rect 113 -428 119 428
rect 73 -440 119 -428
rect 169 428 215 440
rect 169 -428 175 428
rect 209 -428 215 428
rect 169 -440 215 -428
rect 265 428 311 440
rect 265 -428 271 428
rect 305 -428 311 428
rect 265 -440 311 -428
rect 361 428 407 440
rect 361 -428 367 428
rect 401 -428 407 428
rect 361 -440 407 -428
rect -365 -487 -307 -481
rect -365 -521 -353 -487
rect -319 -521 -307 -487
rect -365 -527 -307 -521
rect -173 -487 -115 -481
rect -173 -521 -161 -487
rect -127 -521 -115 -487
rect -173 -527 -115 -521
rect 19 -487 77 -481
rect 19 -521 31 -487
rect 65 -521 77 -487
rect 19 -527 77 -521
rect 211 -487 269 -481
rect 211 -521 223 -487
rect 257 -521 269 -487
rect 211 -527 269 -521
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -498 -606 498 606
string parameters w 4.4 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
