magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_p >>
rect -91 182 267 288
rect 77 120 99 182
rect 109 120 267 182
rect 41 -48 73 120
rect 77 96 267 120
rect 77 95 99 96
rect 77 59 105 95
rect 109 59 267 96
rect 77 -49 267 59
rect -29 -95 29 -89
rect -29 -129 -17 -95
rect -29 -135 29 -129
<< nwell >>
rect -109 120 109 182
rect -109 96 77 120
rect 99 96 109 120
rect -109 59 109 96
rect -109 -49 77 59
rect 99 -49 109 59
rect -109 -148 109 -49
<< pmos >>
rect -15 -48 15 120
<< pdiff >>
rect -73 87 -15 120
rect -73 53 -61 87
rect -27 53 -15 87
rect -73 19 -15 53
rect -73 -15 -61 19
rect -27 -15 -15 19
rect -73 -48 -15 -15
rect 15 87 73 120
rect 15 53 27 87
rect 61 53 73 87
rect 15 19 73 53
rect 15 -15 27 19
rect 61 -15 73 19
rect 15 -48 73 -15
<< pdiffc >>
rect -61 53 -27 87
rect -61 -15 -27 19
rect 27 53 61 87
rect 27 -15 61 19
<< poly >>
rect -15 120 15 146
rect -15 -79 15 -48
rect -33 -95 33 -79
rect -33 -129 -17 -95
rect 17 -129 33 -95
rect -33 -145 33 -129
<< polycont >>
rect -17 -129 17 -95
<< locali >>
rect -61 89 -27 124
rect -61 19 -27 53
rect -61 -52 -27 -17
rect 27 89 61 124
rect 27 19 61 53
rect 27 -52 61 -17
rect -33 -129 -17 -95
rect 17 -129 33 -95
<< viali >>
rect -61 87 -27 89
rect -61 55 -27 87
rect -61 -15 -27 17
rect -61 -17 -27 -15
rect 27 87 61 89
rect 27 55 61 87
rect 27 -15 61 17
rect 27 -17 61 -15
rect -17 -129 17 -95
<< metal1 >>
rect -67 89 -21 120
rect -67 55 -61 89
rect -27 55 -21 89
rect -67 17 -21 55
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -48 -21 -17
rect 21 89 67 120
rect 21 55 27 89
rect 61 55 67 89
rect 77 59 99 95
rect 21 17 67 55
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -48 67 -17
rect -29 -95 29 -89
rect -29 -129 -17 -95
rect 17 -129 29 -95
rect -29 -135 29 -129
<< end >>
