magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 280 35 712
rect -35 -712 35 -280
<< xpolyres >>
rect -35 -280 35 280
<< viali >>
rect -17 658 17 692
rect -17 586 17 620
rect -17 514 17 548
rect -17 442 17 476
rect -17 370 17 404
rect -17 298 17 332
rect -17 -333 17 -299
rect -17 -405 17 -371
rect -17 -477 17 -443
rect -17 -549 17 -515
rect -17 -621 17 -587
rect -17 -693 17 -659
<< metal1 >>
rect -25 692 25 706
rect -25 658 -17 692
rect 17 658 25 692
rect -25 620 25 658
rect -25 586 -17 620
rect 17 586 25 620
rect -25 548 25 586
rect -25 514 -17 548
rect 17 514 25 548
rect -25 476 25 514
rect -25 442 -17 476
rect 17 442 25 476
rect -25 404 25 442
rect -25 370 -17 404
rect 17 370 25 404
rect -25 332 25 370
rect -25 298 -17 332
rect 17 298 25 332
rect -25 285 25 298
rect -25 -299 25 -285
rect -25 -333 -17 -299
rect 17 -333 25 -299
rect -25 -371 25 -333
rect -25 -405 -17 -371
rect 17 -405 25 -371
rect -25 -443 25 -405
rect -25 -477 -17 -443
rect 17 -477 25 -443
rect -25 -515 25 -477
rect -25 -549 -17 -515
rect 17 -549 25 -515
rect -25 -587 25 -549
rect -25 -621 -17 -587
rect 17 -621 25 -587
rect -25 -659 25 -621
rect -25 -693 -17 -659
rect 17 -693 25 -659
rect -25 -706 25 -693
<< end >>
