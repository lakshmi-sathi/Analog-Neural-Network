magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 292 35 724
rect -35 -724 35 -292
<< ppolyres >>
rect -35 -292 35 292
<< viali >>
rect -17 670 17 704
rect -17 598 17 632
rect -17 526 17 560
rect -17 454 17 488
rect -17 382 17 416
rect -17 310 17 344
rect -17 -345 17 -311
rect -17 -417 17 -383
rect -17 -489 17 -455
rect -17 -561 17 -527
rect -17 -633 17 -599
rect -17 -705 17 -671
<< metal1 >>
rect -25 704 25 718
rect -25 670 -17 704
rect 17 670 25 704
rect -25 632 25 670
rect -25 598 -17 632
rect 17 598 25 632
rect -25 560 25 598
rect -25 526 -17 560
rect 17 526 25 560
rect -25 488 25 526
rect -25 454 -17 488
rect 17 454 25 488
rect -25 416 25 454
rect -25 382 -17 416
rect 17 382 25 416
rect -25 344 25 382
rect -25 310 -17 344
rect 17 310 25 344
rect -25 297 25 310
rect -25 -311 25 -297
rect -25 -345 -17 -311
rect 17 -345 25 -311
rect -25 -383 25 -345
rect -25 -417 -17 -383
rect 17 -417 25 -383
rect -25 -455 25 -417
rect -25 -489 -17 -455
rect 17 -489 25 -455
rect -25 -527 25 -489
rect -25 -561 -17 -527
rect 17 -561 25 -527
rect -25 -599 25 -561
rect -25 -633 -17 -599
rect 17 -633 25 -599
rect -25 -671 25 -633
rect -25 -705 -17 -671
rect 17 -705 25 -671
rect -25 -718 25 -705
<< end >>
