magic
tech sky130A
magscale 1 2
timestamp 1627037519
<< xpolycontact >>
rect -35 688 35 1120
rect -35 -1120 35 -688
<< xpolyres >>
rect -35 -688 35 688
<< viali >>
rect -19 705 19 1102
rect -19 -1102 19 -705
<< metal1 >>
rect -25 1102 25 1114
rect -25 705 -19 1102
rect 19 705 25 1102
rect -25 693 25 705
rect -25 -705 25 -693
rect -25 -1102 -19 -705
rect 19 -1102 25 -705
rect -25 -1114 25 -1102
<< res0p35 >>
rect -37 -690 37 690
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 6.88 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 40.0k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
