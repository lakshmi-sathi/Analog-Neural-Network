magic
tech sky130A
magscale 1 2
timestamp 1627921586
<< xpolycontact >>
rect -35 835 35 1267
rect -35 -1267 35 -835
<< xpolyres >>
rect -35 -835 35 835
<< viali >>
rect -19 852 19 1249
rect -19 -1249 19 -852
<< metal1 >>
rect -25 1249 25 1261
rect -25 852 -19 1249
rect 19 852 25 1249
rect -25 840 25 852
rect -25 -852 25 -840
rect -25 -1249 -19 -852
rect 19 -1249 25 -852
rect -25 -1261 25 -1249
<< res0p35 >>
rect -37 -837 37 837
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 8.35 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 48.4k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
