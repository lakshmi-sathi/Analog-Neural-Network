magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< nwell >>
rect 124 792 188 1230
rect 316 792 380 1230
rect 508 792 572 1230
rect 700 792 764 1230
rect 892 792 956 1230
rect 1084 792 1148 1230
rect 1276 792 1340 1230
rect 1468 792 1532 1230
rect 1660 792 1724 1230
rect 124 114 188 552
rect 316 114 380 552
rect 508 114 572 552
rect 700 114 764 552
rect 892 114 956 552
rect 1084 114 1148 552
rect 1276 114 1340 552
rect 1468 114 1532 552
rect 1660 114 1724 552
<< pdiff >>
rect 124 1199 188 1230
rect 124 1165 140 1199
rect 174 1165 188 1199
rect 124 1131 188 1165
rect 124 1097 140 1131
rect 174 1097 188 1131
rect 124 1063 188 1097
rect 124 1029 140 1063
rect 174 1029 188 1063
rect 124 995 188 1029
rect 124 961 140 995
rect 174 961 188 995
rect 124 927 188 961
rect 124 893 140 927
rect 174 893 188 927
rect 124 859 188 893
rect 124 825 140 859
rect 174 825 188 859
rect 124 792 188 825
rect 316 1199 380 1230
rect 316 1165 332 1199
rect 366 1165 380 1199
rect 316 1131 380 1165
rect 316 1097 332 1131
rect 366 1097 380 1131
rect 316 1063 380 1097
rect 316 1029 332 1063
rect 366 1029 380 1063
rect 316 995 380 1029
rect 316 961 332 995
rect 366 961 380 995
rect 316 927 380 961
rect 316 893 332 927
rect 366 893 380 927
rect 316 859 380 893
rect 316 825 332 859
rect 366 825 380 859
rect 316 792 380 825
rect 508 1199 572 1230
rect 508 1165 524 1199
rect 558 1165 572 1199
rect 508 1131 572 1165
rect 508 1097 524 1131
rect 558 1097 572 1131
rect 508 1063 572 1097
rect 508 1029 524 1063
rect 558 1029 572 1063
rect 508 995 572 1029
rect 508 961 524 995
rect 558 961 572 995
rect 508 927 572 961
rect 508 893 524 927
rect 558 893 572 927
rect 508 859 572 893
rect 508 825 524 859
rect 558 825 572 859
rect 508 792 572 825
rect 700 1199 764 1230
rect 700 1165 716 1199
rect 750 1165 764 1199
rect 700 1131 764 1165
rect 700 1097 716 1131
rect 750 1097 764 1131
rect 700 1063 764 1097
rect 700 1029 716 1063
rect 750 1029 764 1063
rect 700 995 764 1029
rect 700 961 716 995
rect 750 961 764 995
rect 700 927 764 961
rect 700 893 716 927
rect 750 893 764 927
rect 700 859 764 893
rect 700 825 716 859
rect 750 825 764 859
rect 700 792 764 825
rect 892 1199 956 1230
rect 892 1165 908 1199
rect 942 1165 956 1199
rect 892 1131 956 1165
rect 892 1097 908 1131
rect 942 1097 956 1131
rect 892 1063 956 1097
rect 892 1029 908 1063
rect 942 1029 956 1063
rect 892 995 956 1029
rect 892 961 908 995
rect 942 961 956 995
rect 892 927 956 961
rect 892 893 908 927
rect 942 893 956 927
rect 892 859 956 893
rect 892 825 908 859
rect 942 825 956 859
rect 892 792 956 825
rect 1084 1199 1148 1230
rect 1084 1165 1100 1199
rect 1134 1165 1148 1199
rect 1084 1131 1148 1165
rect 1084 1097 1100 1131
rect 1134 1097 1148 1131
rect 1084 1063 1148 1097
rect 1084 1029 1100 1063
rect 1134 1029 1148 1063
rect 1084 995 1148 1029
rect 1084 961 1100 995
rect 1134 961 1148 995
rect 1084 927 1148 961
rect 1084 893 1100 927
rect 1134 893 1148 927
rect 1084 859 1148 893
rect 1084 825 1100 859
rect 1134 825 1148 859
rect 1084 792 1148 825
rect 1276 1199 1340 1230
rect 1276 1165 1292 1199
rect 1326 1165 1340 1199
rect 1276 1131 1340 1165
rect 1276 1097 1292 1131
rect 1326 1097 1340 1131
rect 1276 1063 1340 1097
rect 1276 1029 1292 1063
rect 1326 1029 1340 1063
rect 1276 995 1340 1029
rect 1276 961 1292 995
rect 1326 961 1340 995
rect 1276 927 1340 961
rect 1276 893 1292 927
rect 1326 893 1340 927
rect 1276 859 1340 893
rect 1276 825 1292 859
rect 1326 825 1340 859
rect 1276 792 1340 825
rect 1468 1199 1532 1230
rect 1468 1165 1484 1199
rect 1518 1165 1532 1199
rect 1468 1131 1532 1165
rect 1468 1097 1484 1131
rect 1518 1097 1532 1131
rect 1468 1063 1532 1097
rect 1468 1029 1484 1063
rect 1518 1029 1532 1063
rect 1468 995 1532 1029
rect 1468 961 1484 995
rect 1518 961 1532 995
rect 1468 927 1532 961
rect 1468 893 1484 927
rect 1518 893 1532 927
rect 1468 859 1532 893
rect 1468 825 1484 859
rect 1518 825 1532 859
rect 1468 792 1532 825
rect 1660 1199 1724 1230
rect 1660 1165 1676 1199
rect 1710 1165 1724 1199
rect 1660 1131 1724 1165
rect 1660 1097 1676 1131
rect 1710 1097 1724 1131
rect 1660 1063 1724 1097
rect 1660 1029 1676 1063
rect 1710 1029 1724 1063
rect 1660 995 1724 1029
rect 1660 961 1676 995
rect 1710 961 1724 995
rect 1660 927 1724 961
rect 1660 893 1676 927
rect 1710 893 1724 927
rect 1660 859 1724 893
rect 1660 825 1676 859
rect 1710 825 1724 859
rect 1660 792 1724 825
rect 124 521 188 552
rect 124 487 140 521
rect 174 487 188 521
rect 124 453 188 487
rect 124 419 140 453
rect 174 419 188 453
rect 124 385 188 419
rect 124 351 140 385
rect 174 351 188 385
rect 124 317 188 351
rect 124 283 140 317
rect 174 283 188 317
rect 124 249 188 283
rect 124 215 140 249
rect 174 215 188 249
rect 124 181 188 215
rect 124 147 140 181
rect 174 147 188 181
rect 124 114 188 147
rect 316 521 380 552
rect 316 487 332 521
rect 366 487 380 521
rect 316 453 380 487
rect 316 419 332 453
rect 366 419 380 453
rect 316 385 380 419
rect 316 351 332 385
rect 366 351 380 385
rect 316 317 380 351
rect 316 283 332 317
rect 366 283 380 317
rect 316 249 380 283
rect 316 215 332 249
rect 366 215 380 249
rect 316 181 380 215
rect 316 147 332 181
rect 366 147 380 181
rect 316 114 380 147
rect 508 521 572 552
rect 508 487 524 521
rect 558 487 572 521
rect 508 453 572 487
rect 508 419 524 453
rect 558 419 572 453
rect 508 385 572 419
rect 508 351 524 385
rect 558 351 572 385
rect 508 317 572 351
rect 508 283 524 317
rect 558 283 572 317
rect 508 249 572 283
rect 508 215 524 249
rect 558 215 572 249
rect 508 181 572 215
rect 508 147 524 181
rect 558 147 572 181
rect 508 114 572 147
rect 700 521 764 552
rect 700 487 716 521
rect 750 487 764 521
rect 700 453 764 487
rect 700 419 716 453
rect 750 419 764 453
rect 700 385 764 419
rect 700 351 716 385
rect 750 351 764 385
rect 700 317 764 351
rect 700 283 716 317
rect 750 283 764 317
rect 700 249 764 283
rect 700 215 716 249
rect 750 215 764 249
rect 700 181 764 215
rect 700 147 716 181
rect 750 147 764 181
rect 700 114 764 147
rect 892 521 956 552
rect 892 487 908 521
rect 942 487 956 521
rect 892 453 956 487
rect 892 419 908 453
rect 942 419 956 453
rect 892 385 956 419
rect 892 351 908 385
rect 942 351 956 385
rect 892 317 956 351
rect 892 283 908 317
rect 942 283 956 317
rect 892 249 956 283
rect 892 215 908 249
rect 942 215 956 249
rect 892 181 956 215
rect 892 147 908 181
rect 942 147 956 181
rect 892 114 956 147
rect 1084 521 1148 552
rect 1084 487 1100 521
rect 1134 487 1148 521
rect 1084 453 1148 487
rect 1084 419 1100 453
rect 1134 419 1148 453
rect 1084 385 1148 419
rect 1084 351 1100 385
rect 1134 351 1148 385
rect 1084 317 1148 351
rect 1084 283 1100 317
rect 1134 283 1148 317
rect 1084 249 1148 283
rect 1084 215 1100 249
rect 1134 215 1148 249
rect 1084 181 1148 215
rect 1084 147 1100 181
rect 1134 147 1148 181
rect 1084 114 1148 147
rect 1276 521 1340 552
rect 1276 487 1292 521
rect 1326 487 1340 521
rect 1276 453 1340 487
rect 1276 419 1292 453
rect 1326 419 1340 453
rect 1276 385 1340 419
rect 1276 351 1292 385
rect 1326 351 1340 385
rect 1276 317 1340 351
rect 1276 283 1292 317
rect 1326 283 1340 317
rect 1276 249 1340 283
rect 1276 215 1292 249
rect 1326 215 1340 249
rect 1276 181 1340 215
rect 1276 147 1292 181
rect 1326 147 1340 181
rect 1276 114 1340 147
rect 1468 521 1532 552
rect 1468 487 1484 521
rect 1518 487 1532 521
rect 1468 453 1532 487
rect 1468 419 1484 453
rect 1518 419 1532 453
rect 1468 385 1532 419
rect 1468 351 1484 385
rect 1518 351 1532 385
rect 1468 317 1532 351
rect 1468 283 1484 317
rect 1518 283 1532 317
rect 1468 249 1532 283
rect 1468 215 1484 249
rect 1518 215 1532 249
rect 1468 181 1532 215
rect 1468 147 1484 181
rect 1518 147 1532 181
rect 1468 114 1532 147
rect 1660 521 1724 552
rect 1660 487 1676 521
rect 1710 487 1724 521
rect 1660 453 1724 487
rect 1660 419 1676 453
rect 1710 419 1724 453
rect 1660 385 1724 419
rect 1660 351 1676 385
rect 1710 351 1724 385
rect 1660 317 1724 351
rect 1660 283 1676 317
rect 1710 283 1724 317
rect 1660 249 1724 283
rect 1660 215 1676 249
rect 1710 215 1724 249
rect 1660 181 1724 215
rect 1660 147 1676 181
rect 1710 147 1724 181
rect 1660 114 1724 147
<< pdiffc >>
rect 140 1165 174 1199
rect 140 1097 174 1131
rect 140 1029 174 1063
rect 140 961 174 995
rect 140 893 174 927
rect 140 825 174 859
rect 332 1165 366 1199
rect 332 1097 366 1131
rect 332 1029 366 1063
rect 332 961 366 995
rect 332 893 366 927
rect 332 825 366 859
rect 524 1165 558 1199
rect 524 1097 558 1131
rect 524 1029 558 1063
rect 524 961 558 995
rect 524 893 558 927
rect 524 825 558 859
rect 716 1165 750 1199
rect 716 1097 750 1131
rect 716 1029 750 1063
rect 716 961 750 995
rect 716 893 750 927
rect 716 825 750 859
rect 908 1165 942 1199
rect 908 1097 942 1131
rect 908 1029 942 1063
rect 908 961 942 995
rect 908 893 942 927
rect 908 825 942 859
rect 1100 1165 1134 1199
rect 1100 1097 1134 1131
rect 1100 1029 1134 1063
rect 1100 961 1134 995
rect 1100 893 1134 927
rect 1100 825 1134 859
rect 1292 1165 1326 1199
rect 1292 1097 1326 1131
rect 1292 1029 1326 1063
rect 1292 961 1326 995
rect 1292 893 1326 927
rect 1292 825 1326 859
rect 1484 1165 1518 1199
rect 1484 1097 1518 1131
rect 1484 1029 1518 1063
rect 1484 961 1518 995
rect 1484 893 1518 927
rect 1484 825 1518 859
rect 1676 1165 1710 1199
rect 1676 1097 1710 1131
rect 1676 1029 1710 1063
rect 1676 961 1710 995
rect 1676 893 1710 927
rect 1676 825 1710 859
rect 140 487 174 521
rect 140 419 174 453
rect 140 351 174 385
rect 140 283 174 317
rect 140 215 174 249
rect 140 147 174 181
rect 332 487 366 521
rect 332 419 366 453
rect 332 351 366 385
rect 332 283 366 317
rect 332 215 366 249
rect 332 147 366 181
rect 524 487 558 521
rect 524 419 558 453
rect 524 351 558 385
rect 524 283 558 317
rect 524 215 558 249
rect 524 147 558 181
rect 716 487 750 521
rect 716 419 750 453
rect 716 351 750 385
rect 716 283 750 317
rect 716 215 750 249
rect 716 147 750 181
rect 908 487 942 521
rect 908 419 942 453
rect 908 351 942 385
rect 908 283 942 317
rect 908 215 942 249
rect 908 147 942 181
rect 1100 487 1134 521
rect 1100 419 1134 453
rect 1100 351 1134 385
rect 1100 283 1134 317
rect 1100 215 1134 249
rect 1100 147 1134 181
rect 1292 487 1326 521
rect 1292 419 1326 453
rect 1292 351 1326 385
rect 1292 283 1326 317
rect 1292 215 1326 249
rect 1292 147 1326 181
rect 1484 487 1518 521
rect 1484 419 1518 453
rect 1484 351 1518 385
rect 1484 283 1518 317
rect 1484 215 1518 249
rect 1484 147 1518 181
rect 1676 487 1710 521
rect 1676 419 1710 453
rect 1676 351 1710 385
rect 1676 283 1710 317
rect 1676 215 1710 249
rect 1676 147 1710 181
<< poly >>
rect 1659 1289 1756 1315
rect 1665 1285 1756 1289
rect 1726 1233 1756 1285
rect 1726 59 1756 113
rect 1673 55 1756 59
rect 1663 29 1756 55
rect 1665 -305 1760 -279
rect 1675 -309 1760 -305
rect 1730 -340 1760 -309
rect 1730 -987 1760 -942
rect 1669 -1017 1760 -987
<< locali >>
rect -72 1522 1920 1538
rect -72 1488 -67 1522
rect -33 1488 5 1522
rect 39 1488 77 1522
rect 111 1488 149 1522
rect 183 1488 221 1522
rect 255 1488 293 1522
rect 327 1488 365 1522
rect 399 1488 437 1522
rect 471 1488 509 1522
rect 543 1488 581 1522
rect 615 1488 653 1522
rect 687 1488 725 1522
rect 759 1488 797 1522
rect 831 1488 869 1522
rect 903 1488 941 1522
rect 975 1488 1013 1522
rect 1047 1488 1085 1522
rect 1119 1488 1157 1522
rect 1191 1488 1229 1522
rect 1263 1488 1301 1522
rect 1335 1488 1373 1522
rect 1407 1488 1445 1522
rect 1479 1488 1517 1522
rect 1551 1488 1589 1522
rect 1623 1488 1661 1522
rect 1695 1488 1733 1522
rect 1767 1488 1805 1522
rect 1839 1488 1877 1522
rect 1911 1488 1920 1522
rect -72 1462 1920 1488
rect -70 1388 1920 1462
rect 140 1209 174 1230
rect 140 1137 174 1165
rect 140 1065 174 1097
rect 140 995 174 1029
rect 140 927 174 959
rect 140 859 174 887
rect 140 792 174 815
rect 332 1209 366 1230
rect 332 1137 366 1165
rect 332 1065 366 1097
rect 332 995 366 1029
rect 332 927 366 959
rect 332 859 366 887
rect 332 792 366 815
rect 524 1209 558 1230
rect 524 1137 558 1165
rect 524 1065 558 1097
rect 524 995 558 1029
rect 524 927 558 959
rect 524 859 558 887
rect 524 792 558 815
rect 716 1209 750 1230
rect 716 1137 750 1165
rect 716 1065 750 1097
rect 716 995 750 1029
rect 716 927 750 959
rect 716 859 750 887
rect 716 792 750 815
rect 908 1209 942 1230
rect 908 1137 942 1165
rect 908 1065 942 1097
rect 908 995 942 1029
rect 908 927 942 959
rect 908 859 942 887
rect 908 792 942 815
rect 1100 1209 1134 1230
rect 1100 1137 1134 1165
rect 1100 1065 1134 1097
rect 1100 995 1134 1029
rect 1100 927 1134 959
rect 1100 859 1134 887
rect 1100 792 1134 815
rect 1292 1209 1326 1230
rect 1292 1137 1326 1165
rect 1292 1065 1326 1097
rect 1292 995 1326 1029
rect 1292 927 1326 959
rect 1292 859 1326 887
rect 1292 792 1326 815
rect 1484 1209 1518 1230
rect 1484 1137 1518 1165
rect 1484 1065 1518 1097
rect 1484 995 1518 1029
rect 1484 927 1518 959
rect 1484 859 1518 887
rect 1484 792 1518 815
rect 1676 1209 1710 1230
rect 1676 1137 1710 1165
rect 1676 1065 1710 1097
rect 1676 995 1710 1029
rect 1676 927 1710 959
rect 1676 859 1710 887
rect 1676 792 1710 815
rect 140 531 174 552
rect 140 459 174 487
rect 140 387 174 419
rect 140 317 174 351
rect 140 249 174 281
rect 140 181 174 209
rect 140 114 174 137
rect 332 531 366 552
rect 332 459 366 487
rect 332 387 366 419
rect 332 317 366 351
rect 332 249 366 281
rect 332 181 366 209
rect 332 114 366 137
rect 524 531 558 552
rect 524 459 558 487
rect 524 387 558 419
rect 524 317 558 351
rect 524 249 558 281
rect 524 181 558 209
rect 524 114 558 137
rect 716 531 750 552
rect 716 459 750 487
rect 716 387 750 419
rect 716 317 750 351
rect 716 249 750 281
rect 716 181 750 209
rect 716 114 750 137
rect 908 531 942 552
rect 908 459 942 487
rect 908 387 942 419
rect 908 317 942 351
rect 908 249 942 281
rect 908 181 942 209
rect 908 114 942 137
rect 1100 531 1134 552
rect 1100 459 1134 487
rect 1100 387 1134 419
rect 1100 317 1134 351
rect 1100 249 1134 281
rect 1100 181 1134 209
rect 1100 114 1134 137
rect 1292 531 1326 552
rect 1292 459 1326 487
rect 1292 387 1326 419
rect 1292 317 1326 351
rect 1292 249 1326 281
rect 1292 181 1326 209
rect 1292 114 1326 137
rect 1484 531 1518 552
rect 1484 459 1518 487
rect 1484 387 1518 419
rect 1484 317 1518 351
rect 1484 249 1518 281
rect 1484 181 1518 209
rect 1484 114 1518 137
rect 1676 531 1710 552
rect 1676 459 1710 487
rect 1676 387 1710 419
rect 1676 317 1710 351
rect 1676 249 1710 281
rect 1676 181 1710 209
rect 1676 114 1710 137
rect -74 -1158 1926 -1094
rect -66 -1181 1926 -1158
rect -66 -1200 -25 -1181
rect -64 -1215 -25 -1200
rect 9 -1215 47 -1181
rect 81 -1215 119 -1181
rect 153 -1215 191 -1181
rect 225 -1215 263 -1181
rect 297 -1215 335 -1181
rect 369 -1215 407 -1181
rect 441 -1215 479 -1181
rect 513 -1215 551 -1181
rect 585 -1215 623 -1181
rect 657 -1215 695 -1181
rect 729 -1215 767 -1181
rect 801 -1215 839 -1181
rect 873 -1215 911 -1181
rect 945 -1215 983 -1181
rect 1017 -1215 1055 -1181
rect 1089 -1215 1127 -1181
rect 1161 -1215 1199 -1181
rect 1233 -1215 1271 -1181
rect 1305 -1215 1343 -1181
rect 1377 -1215 1415 -1181
rect 1449 -1215 1487 -1181
rect 1521 -1215 1559 -1181
rect 1593 -1215 1631 -1181
rect 1665 -1215 1703 -1181
rect 1737 -1215 1775 -1181
rect 1809 -1215 1847 -1181
rect 1881 -1215 1926 -1181
rect -64 -1242 1926 -1215
<< viali >>
rect -67 1488 -33 1522
rect 5 1488 39 1522
rect 77 1488 111 1522
rect 149 1488 183 1522
rect 221 1488 255 1522
rect 293 1488 327 1522
rect 365 1488 399 1522
rect 437 1488 471 1522
rect 509 1488 543 1522
rect 581 1488 615 1522
rect 653 1488 687 1522
rect 725 1488 759 1522
rect 797 1488 831 1522
rect 869 1488 903 1522
rect 941 1488 975 1522
rect 1013 1488 1047 1522
rect 1085 1488 1119 1522
rect 1157 1488 1191 1522
rect 1229 1488 1263 1522
rect 1301 1488 1335 1522
rect 1373 1488 1407 1522
rect 1445 1488 1479 1522
rect 1517 1488 1551 1522
rect 1589 1488 1623 1522
rect 1661 1488 1695 1522
rect 1733 1488 1767 1522
rect 1805 1488 1839 1522
rect 1877 1488 1911 1522
rect 140 1199 174 1209
rect 140 1175 174 1199
rect 140 1131 174 1137
rect 140 1103 174 1131
rect 140 1063 174 1065
rect 140 1031 174 1063
rect 140 961 174 993
rect 140 959 174 961
rect 140 893 174 921
rect 140 887 174 893
rect 140 825 174 849
rect 140 815 174 825
rect 332 1199 366 1209
rect 332 1175 366 1199
rect 332 1131 366 1137
rect 332 1103 366 1131
rect 332 1063 366 1065
rect 332 1031 366 1063
rect 332 961 366 993
rect 332 959 366 961
rect 332 893 366 921
rect 332 887 366 893
rect 332 825 366 849
rect 332 815 366 825
rect 524 1199 558 1209
rect 524 1175 558 1199
rect 524 1131 558 1137
rect 524 1103 558 1131
rect 524 1063 558 1065
rect 524 1031 558 1063
rect 524 961 558 993
rect 524 959 558 961
rect 524 893 558 921
rect 524 887 558 893
rect 524 825 558 849
rect 524 815 558 825
rect 716 1199 750 1209
rect 716 1175 750 1199
rect 716 1131 750 1137
rect 716 1103 750 1131
rect 716 1063 750 1065
rect 716 1031 750 1063
rect 716 961 750 993
rect 716 959 750 961
rect 716 893 750 921
rect 716 887 750 893
rect 716 825 750 849
rect 716 815 750 825
rect 908 1199 942 1209
rect 908 1175 942 1199
rect 908 1131 942 1137
rect 908 1103 942 1131
rect 908 1063 942 1065
rect 908 1031 942 1063
rect 908 961 942 993
rect 908 959 942 961
rect 908 893 942 921
rect 908 887 942 893
rect 908 825 942 849
rect 908 815 942 825
rect 1100 1199 1134 1209
rect 1100 1175 1134 1199
rect 1100 1131 1134 1137
rect 1100 1103 1134 1131
rect 1100 1063 1134 1065
rect 1100 1031 1134 1063
rect 1100 961 1134 993
rect 1100 959 1134 961
rect 1100 893 1134 921
rect 1100 887 1134 893
rect 1100 825 1134 849
rect 1100 815 1134 825
rect 1292 1199 1326 1209
rect 1292 1175 1326 1199
rect 1292 1131 1326 1137
rect 1292 1103 1326 1131
rect 1292 1063 1326 1065
rect 1292 1031 1326 1063
rect 1292 961 1326 993
rect 1292 959 1326 961
rect 1292 893 1326 921
rect 1292 887 1326 893
rect 1292 825 1326 849
rect 1292 815 1326 825
rect 1484 1199 1518 1209
rect 1484 1175 1518 1199
rect 1484 1131 1518 1137
rect 1484 1103 1518 1131
rect 1484 1063 1518 1065
rect 1484 1031 1518 1063
rect 1484 961 1518 993
rect 1484 959 1518 961
rect 1484 893 1518 921
rect 1484 887 1518 893
rect 1484 825 1518 849
rect 1484 815 1518 825
rect 1676 1199 1710 1209
rect 1676 1175 1710 1199
rect 1676 1131 1710 1137
rect 1676 1103 1710 1131
rect 1676 1063 1710 1065
rect 1676 1031 1710 1063
rect 1676 961 1710 993
rect 1676 959 1710 961
rect 1676 893 1710 921
rect 1676 887 1710 893
rect 1676 825 1710 849
rect 1676 815 1710 825
rect 140 521 174 531
rect 140 497 174 521
rect 140 453 174 459
rect 140 425 174 453
rect 140 385 174 387
rect 140 353 174 385
rect 140 283 174 315
rect 140 281 174 283
rect 140 215 174 243
rect 140 209 174 215
rect 140 147 174 171
rect 140 137 174 147
rect 332 521 366 531
rect 332 497 366 521
rect 332 453 366 459
rect 332 425 366 453
rect 332 385 366 387
rect 332 353 366 385
rect 332 283 366 315
rect 332 281 366 283
rect 332 215 366 243
rect 332 209 366 215
rect 332 147 366 171
rect 332 137 366 147
rect 524 521 558 531
rect 524 497 558 521
rect 524 453 558 459
rect 524 425 558 453
rect 524 385 558 387
rect 524 353 558 385
rect 524 283 558 315
rect 524 281 558 283
rect 524 215 558 243
rect 524 209 558 215
rect 524 147 558 171
rect 524 137 558 147
rect 716 521 750 531
rect 716 497 750 521
rect 716 453 750 459
rect 716 425 750 453
rect 716 385 750 387
rect 716 353 750 385
rect 716 283 750 315
rect 716 281 750 283
rect 716 215 750 243
rect 716 209 750 215
rect 716 147 750 171
rect 716 137 750 147
rect 908 521 942 531
rect 908 497 942 521
rect 908 453 942 459
rect 908 425 942 453
rect 908 385 942 387
rect 908 353 942 385
rect 908 283 942 315
rect 908 281 942 283
rect 908 215 942 243
rect 908 209 942 215
rect 908 147 942 171
rect 908 137 942 147
rect 1100 521 1134 531
rect 1100 497 1134 521
rect 1100 453 1134 459
rect 1100 425 1134 453
rect 1100 385 1134 387
rect 1100 353 1134 385
rect 1100 283 1134 315
rect 1100 281 1134 283
rect 1100 215 1134 243
rect 1100 209 1134 215
rect 1100 147 1134 171
rect 1100 137 1134 147
rect 1292 521 1326 531
rect 1292 497 1326 521
rect 1292 453 1326 459
rect 1292 425 1326 453
rect 1292 385 1326 387
rect 1292 353 1326 385
rect 1292 283 1326 315
rect 1292 281 1326 283
rect 1292 215 1326 243
rect 1292 209 1326 215
rect 1292 147 1326 171
rect 1292 137 1326 147
rect 1484 521 1518 531
rect 1484 497 1518 521
rect 1484 453 1518 459
rect 1484 425 1518 453
rect 1484 385 1518 387
rect 1484 353 1518 385
rect 1484 283 1518 315
rect 1484 281 1518 283
rect 1484 215 1518 243
rect 1484 209 1518 215
rect 1484 147 1518 171
rect 1484 137 1518 147
rect 1676 521 1710 531
rect 1676 497 1710 521
rect 1676 453 1710 459
rect 1676 425 1710 453
rect 1676 385 1710 387
rect 1676 353 1710 385
rect 1676 283 1710 315
rect 1676 281 1710 283
rect 1676 215 1710 243
rect 1676 209 1710 215
rect 1676 147 1710 171
rect 1676 137 1710 147
rect -25 -1215 9 -1181
rect 47 -1215 81 -1181
rect 119 -1215 153 -1181
rect 191 -1215 225 -1181
rect 263 -1215 297 -1181
rect 335 -1215 369 -1181
rect 407 -1215 441 -1181
rect 479 -1215 513 -1181
rect 551 -1215 585 -1181
rect 623 -1215 657 -1181
rect 695 -1215 729 -1181
rect 767 -1215 801 -1181
rect 839 -1215 873 -1181
rect 911 -1215 945 -1181
rect 983 -1215 1017 -1181
rect 1055 -1215 1089 -1181
rect 1127 -1215 1161 -1181
rect 1199 -1215 1233 -1181
rect 1271 -1215 1305 -1181
rect 1343 -1215 1377 -1181
rect 1415 -1215 1449 -1181
rect 1487 -1215 1521 -1181
rect 1559 -1215 1593 -1181
rect 1631 -1215 1665 -1181
rect 1703 -1215 1737 -1181
rect 1775 -1215 1809 -1181
rect 1847 -1215 1881 -1181
<< metal1 >>
rect -84 1536 1924 1554
rect -84 1522 -66 1536
rect -84 1488 -67 1522
rect -84 1484 -66 1488
rect -14 1484 -2 1536
rect 50 1484 62 1536
rect 114 1484 126 1536
rect 178 1522 190 1536
rect 242 1522 254 1536
rect 306 1522 318 1536
rect 370 1522 382 1536
rect 434 1522 446 1536
rect 498 1522 510 1536
rect 183 1488 190 1522
rect 434 1488 437 1522
rect 498 1488 509 1522
rect 178 1484 190 1488
rect 242 1484 254 1488
rect 306 1484 318 1488
rect 370 1484 382 1488
rect 434 1484 446 1488
rect 498 1484 510 1488
rect 562 1484 574 1536
rect 626 1484 638 1536
rect 690 1484 702 1536
rect 754 1522 766 1536
rect 818 1522 830 1536
rect 882 1522 894 1536
rect 946 1522 958 1536
rect 1010 1522 1022 1536
rect 1074 1522 1086 1536
rect 759 1488 766 1522
rect 1010 1488 1013 1522
rect 1074 1488 1085 1522
rect 754 1484 766 1488
rect 818 1484 830 1488
rect 882 1484 894 1488
rect 946 1484 958 1488
rect 1010 1484 1022 1488
rect 1074 1484 1086 1488
rect 1138 1484 1150 1536
rect 1202 1484 1214 1536
rect 1266 1484 1278 1536
rect 1330 1522 1342 1536
rect 1394 1522 1406 1536
rect 1458 1522 1470 1536
rect 1522 1522 1534 1536
rect 1586 1522 1598 1536
rect 1650 1522 1662 1536
rect 1335 1488 1342 1522
rect 1586 1488 1589 1522
rect 1650 1488 1661 1522
rect 1330 1484 1342 1488
rect 1394 1484 1406 1488
rect 1458 1484 1470 1488
rect 1522 1484 1534 1488
rect 1586 1484 1598 1488
rect 1650 1484 1662 1488
rect 1714 1484 1726 1536
rect 1778 1484 1790 1536
rect 1842 1484 1854 1536
rect 1906 1522 1924 1536
rect 1911 1488 1924 1522
rect 1906 1484 1924 1488
rect -84 1464 1924 1484
rect 78 1274 1676 1322
rect 30 1195 94 1226
rect 30 1143 36 1195
rect 88 1143 94 1195
rect 30 1131 94 1143
rect 30 1079 36 1131
rect 88 1079 94 1131
rect 30 1067 94 1079
rect 30 1015 36 1067
rect 88 1015 94 1067
rect 30 1003 94 1015
rect 30 951 36 1003
rect 88 951 94 1003
rect 30 939 94 951
rect 30 887 36 939
rect 88 887 94 939
rect 30 875 94 887
rect 30 823 36 875
rect 88 823 94 875
rect 30 792 94 823
rect 124 1209 188 1230
rect 124 1197 140 1209
rect 174 1197 188 1209
rect 124 1145 130 1197
rect 182 1145 188 1197
rect 124 1137 188 1145
rect 124 1133 140 1137
rect 174 1133 188 1137
rect 124 1081 130 1133
rect 182 1081 188 1133
rect 124 1069 188 1081
rect 124 1017 130 1069
rect 182 1017 188 1069
rect 124 1005 188 1017
rect 124 953 130 1005
rect 182 953 188 1005
rect 124 941 188 953
rect 124 889 130 941
rect 182 889 188 941
rect 124 887 140 889
rect 174 887 188 889
rect 124 877 188 887
rect 124 825 130 877
rect 182 825 188 877
rect 124 815 140 825
rect 174 815 188 825
rect 124 792 188 815
rect 222 1195 286 1226
rect 222 1143 228 1195
rect 280 1143 286 1195
rect 222 1131 286 1143
rect 222 1079 228 1131
rect 280 1079 286 1131
rect 222 1067 286 1079
rect 222 1015 228 1067
rect 280 1015 286 1067
rect 222 1003 286 1015
rect 222 951 228 1003
rect 280 951 286 1003
rect 222 939 286 951
rect 222 887 228 939
rect 280 887 286 939
rect 222 875 286 887
rect 222 823 228 875
rect 280 823 286 875
rect 222 792 286 823
rect 316 1209 380 1230
rect 316 1197 332 1209
rect 366 1197 380 1209
rect 316 1145 322 1197
rect 374 1145 380 1197
rect 316 1137 380 1145
rect 316 1133 332 1137
rect 366 1133 380 1137
rect 316 1081 322 1133
rect 374 1081 380 1133
rect 316 1069 380 1081
rect 316 1017 322 1069
rect 374 1017 380 1069
rect 316 1005 380 1017
rect 316 953 322 1005
rect 374 953 380 1005
rect 316 941 380 953
rect 316 889 322 941
rect 374 889 380 941
rect 316 887 332 889
rect 366 887 380 889
rect 316 877 380 887
rect 316 825 322 877
rect 374 825 380 877
rect 316 815 332 825
rect 366 815 380 825
rect 316 792 380 815
rect 414 1195 478 1226
rect 414 1143 420 1195
rect 472 1143 478 1195
rect 414 1131 478 1143
rect 414 1079 420 1131
rect 472 1079 478 1131
rect 414 1067 478 1079
rect 414 1015 420 1067
rect 472 1015 478 1067
rect 414 1003 478 1015
rect 414 951 420 1003
rect 472 951 478 1003
rect 414 939 478 951
rect 414 887 420 939
rect 472 887 478 939
rect 414 875 478 887
rect 414 823 420 875
rect 472 823 478 875
rect 414 792 478 823
rect 508 1209 572 1230
rect 508 1197 524 1209
rect 558 1197 572 1209
rect 508 1145 514 1197
rect 566 1145 572 1197
rect 508 1137 572 1145
rect 508 1133 524 1137
rect 558 1133 572 1137
rect 508 1081 514 1133
rect 566 1081 572 1133
rect 508 1069 572 1081
rect 508 1017 514 1069
rect 566 1017 572 1069
rect 508 1005 572 1017
rect 508 953 514 1005
rect 566 953 572 1005
rect 508 941 572 953
rect 508 889 514 941
rect 566 889 572 941
rect 508 887 524 889
rect 558 887 572 889
rect 508 877 572 887
rect 508 825 514 877
rect 566 825 572 877
rect 508 815 524 825
rect 558 815 572 825
rect 508 792 572 815
rect 606 1195 670 1226
rect 606 1143 612 1195
rect 664 1143 670 1195
rect 606 1131 670 1143
rect 606 1079 612 1131
rect 664 1079 670 1131
rect 606 1067 670 1079
rect 606 1015 612 1067
rect 664 1015 670 1067
rect 606 1003 670 1015
rect 606 951 612 1003
rect 664 951 670 1003
rect 606 939 670 951
rect 606 887 612 939
rect 664 887 670 939
rect 606 875 670 887
rect 606 823 612 875
rect 664 823 670 875
rect 606 792 670 823
rect 700 1209 764 1230
rect 700 1197 716 1209
rect 750 1197 764 1209
rect 700 1145 706 1197
rect 758 1145 764 1197
rect 700 1137 764 1145
rect 700 1133 716 1137
rect 750 1133 764 1137
rect 700 1081 706 1133
rect 758 1081 764 1133
rect 700 1069 764 1081
rect 700 1017 706 1069
rect 758 1017 764 1069
rect 700 1005 764 1017
rect 700 953 706 1005
rect 758 953 764 1005
rect 700 941 764 953
rect 700 889 706 941
rect 758 889 764 941
rect 700 887 716 889
rect 750 887 764 889
rect 700 877 764 887
rect 700 825 706 877
rect 758 825 764 877
rect 700 815 716 825
rect 750 815 764 825
rect 700 792 764 815
rect 798 1195 862 1226
rect 798 1143 804 1195
rect 856 1143 862 1195
rect 798 1131 862 1143
rect 798 1079 804 1131
rect 856 1079 862 1131
rect 798 1067 862 1079
rect 798 1015 804 1067
rect 856 1015 862 1067
rect 798 1003 862 1015
rect 798 951 804 1003
rect 856 951 862 1003
rect 798 939 862 951
rect 798 887 804 939
rect 856 887 862 939
rect 798 875 862 887
rect 798 823 804 875
rect 856 823 862 875
rect 798 792 862 823
rect 892 1209 956 1230
rect 892 1197 908 1209
rect 942 1197 956 1209
rect 892 1145 898 1197
rect 950 1145 956 1197
rect 892 1137 956 1145
rect 892 1133 908 1137
rect 942 1133 956 1137
rect 892 1081 898 1133
rect 950 1081 956 1133
rect 892 1069 956 1081
rect 892 1017 898 1069
rect 950 1017 956 1069
rect 892 1005 956 1017
rect 892 953 898 1005
rect 950 953 956 1005
rect 892 941 956 953
rect 892 889 898 941
rect 950 889 956 941
rect 892 887 908 889
rect 942 887 956 889
rect 892 877 956 887
rect 892 825 898 877
rect 950 825 956 877
rect 892 815 908 825
rect 942 815 956 825
rect 892 792 956 815
rect 990 1195 1054 1226
rect 990 1143 996 1195
rect 1048 1143 1054 1195
rect 990 1131 1054 1143
rect 990 1079 996 1131
rect 1048 1079 1054 1131
rect 990 1067 1054 1079
rect 990 1015 996 1067
rect 1048 1015 1054 1067
rect 990 1003 1054 1015
rect 990 951 996 1003
rect 1048 951 1054 1003
rect 990 939 1054 951
rect 990 887 996 939
rect 1048 887 1054 939
rect 990 875 1054 887
rect 990 823 996 875
rect 1048 823 1054 875
rect 990 792 1054 823
rect 1084 1209 1148 1230
rect 1084 1197 1100 1209
rect 1134 1197 1148 1209
rect 1084 1145 1090 1197
rect 1142 1145 1148 1197
rect 1084 1137 1148 1145
rect 1084 1133 1100 1137
rect 1134 1133 1148 1137
rect 1084 1081 1090 1133
rect 1142 1081 1148 1133
rect 1084 1069 1148 1081
rect 1084 1017 1090 1069
rect 1142 1017 1148 1069
rect 1084 1005 1148 1017
rect 1084 953 1090 1005
rect 1142 953 1148 1005
rect 1084 941 1148 953
rect 1084 889 1090 941
rect 1142 889 1148 941
rect 1084 887 1100 889
rect 1134 887 1148 889
rect 1084 877 1148 887
rect 1084 825 1090 877
rect 1142 825 1148 877
rect 1084 815 1100 825
rect 1134 815 1148 825
rect 1084 792 1148 815
rect 1182 1195 1246 1226
rect 1182 1143 1188 1195
rect 1240 1143 1246 1195
rect 1182 1131 1246 1143
rect 1182 1079 1188 1131
rect 1240 1079 1246 1131
rect 1182 1067 1246 1079
rect 1182 1015 1188 1067
rect 1240 1015 1246 1067
rect 1182 1003 1246 1015
rect 1182 951 1188 1003
rect 1240 951 1246 1003
rect 1182 939 1246 951
rect 1182 887 1188 939
rect 1240 887 1246 939
rect 1182 875 1246 887
rect 1182 823 1188 875
rect 1240 823 1246 875
rect 1182 792 1246 823
rect 1276 1209 1340 1230
rect 1276 1197 1292 1209
rect 1326 1197 1340 1209
rect 1276 1145 1282 1197
rect 1334 1145 1340 1197
rect 1276 1137 1340 1145
rect 1276 1133 1292 1137
rect 1326 1133 1340 1137
rect 1276 1081 1282 1133
rect 1334 1081 1340 1133
rect 1276 1069 1340 1081
rect 1276 1017 1282 1069
rect 1334 1017 1340 1069
rect 1276 1005 1340 1017
rect 1276 953 1282 1005
rect 1334 953 1340 1005
rect 1276 941 1340 953
rect 1276 889 1282 941
rect 1334 889 1340 941
rect 1276 887 1292 889
rect 1326 887 1340 889
rect 1276 877 1340 887
rect 1276 825 1282 877
rect 1334 825 1340 877
rect 1276 815 1292 825
rect 1326 815 1340 825
rect 1276 792 1340 815
rect 1374 1195 1438 1226
rect 1374 1143 1380 1195
rect 1432 1143 1438 1195
rect 1374 1131 1438 1143
rect 1374 1079 1380 1131
rect 1432 1079 1438 1131
rect 1374 1067 1438 1079
rect 1374 1015 1380 1067
rect 1432 1015 1438 1067
rect 1374 1003 1438 1015
rect 1374 951 1380 1003
rect 1432 951 1438 1003
rect 1374 939 1438 951
rect 1374 887 1380 939
rect 1432 887 1438 939
rect 1374 875 1438 887
rect 1374 823 1380 875
rect 1432 823 1438 875
rect 1374 792 1438 823
rect 1468 1209 1532 1230
rect 1468 1197 1484 1209
rect 1518 1197 1532 1209
rect 1468 1145 1474 1197
rect 1526 1145 1532 1197
rect 1468 1137 1532 1145
rect 1468 1133 1484 1137
rect 1518 1133 1532 1137
rect 1468 1081 1474 1133
rect 1526 1081 1532 1133
rect 1468 1069 1532 1081
rect 1468 1017 1474 1069
rect 1526 1017 1532 1069
rect 1468 1005 1532 1017
rect 1468 953 1474 1005
rect 1526 953 1532 1005
rect 1468 941 1532 953
rect 1468 889 1474 941
rect 1526 889 1532 941
rect 1468 887 1484 889
rect 1518 887 1532 889
rect 1468 877 1532 887
rect 1468 825 1474 877
rect 1526 825 1532 877
rect 1468 815 1484 825
rect 1518 815 1532 825
rect 1468 792 1532 815
rect 1566 1195 1630 1226
rect 1566 1143 1572 1195
rect 1624 1143 1630 1195
rect 1566 1131 1630 1143
rect 1566 1079 1572 1131
rect 1624 1079 1630 1131
rect 1566 1067 1630 1079
rect 1566 1015 1572 1067
rect 1624 1015 1630 1067
rect 1566 1003 1630 1015
rect 1566 951 1572 1003
rect 1624 951 1630 1003
rect 1566 939 1630 951
rect 1566 887 1572 939
rect 1624 887 1630 939
rect 1566 875 1630 887
rect 1566 823 1572 875
rect 1624 823 1630 875
rect 1566 792 1630 823
rect 1660 1209 1724 1230
rect 1660 1197 1676 1209
rect 1710 1197 1724 1209
rect 1660 1145 1666 1197
rect 1718 1145 1724 1197
rect 1660 1137 1724 1145
rect 1660 1133 1676 1137
rect 1710 1133 1724 1137
rect 1660 1081 1666 1133
rect 1718 1081 1724 1133
rect 1660 1069 1724 1081
rect 1660 1017 1666 1069
rect 1718 1017 1724 1069
rect 1660 1005 1724 1017
rect 1660 953 1666 1005
rect 1718 953 1724 1005
rect 1660 941 1724 953
rect 1660 889 1666 941
rect 1718 889 1724 941
rect 1660 887 1676 889
rect 1710 887 1724 889
rect 1660 877 1724 887
rect 1660 825 1666 877
rect 1718 825 1724 877
rect 1660 815 1676 825
rect 1710 815 1724 825
rect 1660 792 1724 815
rect 1758 1195 1822 1226
rect 1758 1143 1764 1195
rect 1816 1143 1822 1195
rect 1758 1131 1822 1143
rect 1758 1079 1764 1131
rect 1816 1079 1822 1131
rect 1758 1067 1822 1079
rect 1758 1015 1764 1067
rect 1816 1015 1822 1067
rect 1758 1003 1822 1015
rect 1758 951 1764 1003
rect 1816 951 1822 1003
rect 1758 939 1822 951
rect 1758 887 1764 939
rect 1816 887 1822 939
rect 1758 875 1822 887
rect 1758 823 1764 875
rect 1816 823 1822 875
rect 1758 792 1822 823
rect -166 596 1772 752
rect -166 -564 -10 596
rect 30 517 94 548
rect 30 465 36 517
rect 88 465 94 517
rect 30 453 94 465
rect 30 401 36 453
rect 88 401 94 453
rect 30 389 94 401
rect 30 337 36 389
rect 88 337 94 389
rect 30 325 94 337
rect 30 273 36 325
rect 88 273 94 325
rect 30 261 94 273
rect 30 209 36 261
rect 88 209 94 261
rect 30 197 94 209
rect 30 145 36 197
rect 88 145 94 197
rect 30 114 94 145
rect 124 531 188 552
rect 124 519 140 531
rect 174 519 188 531
rect 124 467 130 519
rect 182 467 188 519
rect 124 459 188 467
rect 124 455 140 459
rect 174 455 188 459
rect 124 403 130 455
rect 182 403 188 455
rect 124 391 188 403
rect 124 339 130 391
rect 182 339 188 391
rect 124 327 188 339
rect 124 275 130 327
rect 182 275 188 327
rect 124 263 188 275
rect 124 211 130 263
rect 182 211 188 263
rect 124 209 140 211
rect 174 209 188 211
rect 124 199 188 209
rect 124 147 130 199
rect 182 147 188 199
rect 124 137 140 147
rect 174 137 188 147
rect 124 114 188 137
rect 222 517 286 548
rect 222 465 228 517
rect 280 465 286 517
rect 222 453 286 465
rect 222 401 228 453
rect 280 401 286 453
rect 222 389 286 401
rect 222 337 228 389
rect 280 337 286 389
rect 222 325 286 337
rect 222 273 228 325
rect 280 273 286 325
rect 222 261 286 273
rect 222 209 228 261
rect 280 209 286 261
rect 222 197 286 209
rect 222 145 228 197
rect 280 145 286 197
rect 222 114 286 145
rect 316 531 380 552
rect 316 519 332 531
rect 366 519 380 531
rect 316 467 322 519
rect 374 467 380 519
rect 316 459 380 467
rect 316 455 332 459
rect 366 455 380 459
rect 316 403 322 455
rect 374 403 380 455
rect 316 391 380 403
rect 316 339 322 391
rect 374 339 380 391
rect 316 327 380 339
rect 316 275 322 327
rect 374 275 380 327
rect 316 263 380 275
rect 316 211 322 263
rect 374 211 380 263
rect 316 209 332 211
rect 366 209 380 211
rect 316 199 380 209
rect 316 147 322 199
rect 374 147 380 199
rect 316 137 332 147
rect 366 137 380 147
rect 316 114 380 137
rect 414 517 478 548
rect 414 465 420 517
rect 472 465 478 517
rect 414 453 478 465
rect 414 401 420 453
rect 472 401 478 453
rect 414 389 478 401
rect 414 337 420 389
rect 472 337 478 389
rect 414 325 478 337
rect 414 273 420 325
rect 472 273 478 325
rect 414 261 478 273
rect 414 209 420 261
rect 472 209 478 261
rect 414 197 478 209
rect 414 145 420 197
rect 472 145 478 197
rect 414 114 478 145
rect 508 531 572 552
rect 508 519 524 531
rect 558 519 572 531
rect 508 467 514 519
rect 566 467 572 519
rect 508 459 572 467
rect 508 455 524 459
rect 558 455 572 459
rect 508 403 514 455
rect 566 403 572 455
rect 508 391 572 403
rect 508 339 514 391
rect 566 339 572 391
rect 508 327 572 339
rect 508 275 514 327
rect 566 275 572 327
rect 508 263 572 275
rect 508 211 514 263
rect 566 211 572 263
rect 508 209 524 211
rect 558 209 572 211
rect 508 199 572 209
rect 508 147 514 199
rect 566 147 572 199
rect 508 137 524 147
rect 558 137 572 147
rect 508 114 572 137
rect 606 517 670 548
rect 606 465 612 517
rect 664 465 670 517
rect 606 453 670 465
rect 606 401 612 453
rect 664 401 670 453
rect 606 389 670 401
rect 606 337 612 389
rect 664 337 670 389
rect 606 325 670 337
rect 606 273 612 325
rect 664 273 670 325
rect 606 261 670 273
rect 606 209 612 261
rect 664 209 670 261
rect 606 197 670 209
rect 606 145 612 197
rect 664 145 670 197
rect 606 114 670 145
rect 700 531 764 552
rect 700 519 716 531
rect 750 519 764 531
rect 700 467 706 519
rect 758 467 764 519
rect 700 459 764 467
rect 700 455 716 459
rect 750 455 764 459
rect 700 403 706 455
rect 758 403 764 455
rect 700 391 764 403
rect 700 339 706 391
rect 758 339 764 391
rect 700 327 764 339
rect 700 275 706 327
rect 758 275 764 327
rect 700 263 764 275
rect 700 211 706 263
rect 758 211 764 263
rect 700 209 716 211
rect 750 209 764 211
rect 700 199 764 209
rect 700 147 706 199
rect 758 147 764 199
rect 700 137 716 147
rect 750 137 764 147
rect 700 114 764 137
rect 798 517 862 548
rect 798 465 804 517
rect 856 465 862 517
rect 798 453 862 465
rect 798 401 804 453
rect 856 401 862 453
rect 798 389 862 401
rect 798 337 804 389
rect 856 337 862 389
rect 798 325 862 337
rect 798 273 804 325
rect 856 273 862 325
rect 798 261 862 273
rect 798 209 804 261
rect 856 209 862 261
rect 798 197 862 209
rect 798 145 804 197
rect 856 145 862 197
rect 798 114 862 145
rect 892 531 956 552
rect 892 519 908 531
rect 942 519 956 531
rect 892 467 898 519
rect 950 467 956 519
rect 892 459 956 467
rect 892 455 908 459
rect 942 455 956 459
rect 892 403 898 455
rect 950 403 956 455
rect 892 391 956 403
rect 892 339 898 391
rect 950 339 956 391
rect 892 327 956 339
rect 892 275 898 327
rect 950 275 956 327
rect 892 263 956 275
rect 892 211 898 263
rect 950 211 956 263
rect 892 209 908 211
rect 942 209 956 211
rect 892 199 956 209
rect 892 147 898 199
rect 950 147 956 199
rect 892 137 908 147
rect 942 137 956 147
rect 892 114 956 137
rect 990 517 1054 548
rect 990 465 996 517
rect 1048 465 1054 517
rect 990 453 1054 465
rect 990 401 996 453
rect 1048 401 1054 453
rect 990 389 1054 401
rect 990 337 996 389
rect 1048 337 1054 389
rect 990 325 1054 337
rect 990 273 996 325
rect 1048 273 1054 325
rect 990 261 1054 273
rect 990 209 996 261
rect 1048 209 1054 261
rect 990 197 1054 209
rect 990 145 996 197
rect 1048 145 1054 197
rect 990 114 1054 145
rect 1084 531 1148 552
rect 1084 519 1100 531
rect 1134 519 1148 531
rect 1084 467 1090 519
rect 1142 467 1148 519
rect 1084 459 1148 467
rect 1084 455 1100 459
rect 1134 455 1148 459
rect 1084 403 1090 455
rect 1142 403 1148 455
rect 1084 391 1148 403
rect 1084 339 1090 391
rect 1142 339 1148 391
rect 1084 327 1148 339
rect 1084 275 1090 327
rect 1142 275 1148 327
rect 1084 263 1148 275
rect 1084 211 1090 263
rect 1142 211 1148 263
rect 1084 209 1100 211
rect 1134 209 1148 211
rect 1084 199 1148 209
rect 1084 147 1090 199
rect 1142 147 1148 199
rect 1084 137 1100 147
rect 1134 137 1148 147
rect 1084 114 1148 137
rect 1182 517 1246 548
rect 1182 465 1188 517
rect 1240 465 1246 517
rect 1182 453 1246 465
rect 1182 401 1188 453
rect 1240 401 1246 453
rect 1182 389 1246 401
rect 1182 337 1188 389
rect 1240 337 1246 389
rect 1182 325 1246 337
rect 1182 273 1188 325
rect 1240 273 1246 325
rect 1182 261 1246 273
rect 1182 209 1188 261
rect 1240 209 1246 261
rect 1182 197 1246 209
rect 1182 145 1188 197
rect 1240 145 1246 197
rect 1182 114 1246 145
rect 1276 531 1340 552
rect 1276 519 1292 531
rect 1326 519 1340 531
rect 1276 467 1282 519
rect 1334 467 1340 519
rect 1276 459 1340 467
rect 1276 455 1292 459
rect 1326 455 1340 459
rect 1276 403 1282 455
rect 1334 403 1340 455
rect 1276 391 1340 403
rect 1276 339 1282 391
rect 1334 339 1340 391
rect 1276 327 1340 339
rect 1276 275 1282 327
rect 1334 275 1340 327
rect 1276 263 1340 275
rect 1276 211 1282 263
rect 1334 211 1340 263
rect 1276 209 1292 211
rect 1326 209 1340 211
rect 1276 199 1340 209
rect 1276 147 1282 199
rect 1334 147 1340 199
rect 1276 137 1292 147
rect 1326 137 1340 147
rect 1276 114 1340 137
rect 1374 517 1438 548
rect 1374 465 1380 517
rect 1432 465 1438 517
rect 1374 453 1438 465
rect 1374 401 1380 453
rect 1432 401 1438 453
rect 1374 389 1438 401
rect 1374 337 1380 389
rect 1432 337 1438 389
rect 1374 325 1438 337
rect 1374 273 1380 325
rect 1432 273 1438 325
rect 1374 261 1438 273
rect 1374 209 1380 261
rect 1432 209 1438 261
rect 1374 197 1438 209
rect 1374 145 1380 197
rect 1432 145 1438 197
rect 1374 114 1438 145
rect 1468 531 1532 552
rect 1468 519 1484 531
rect 1518 519 1532 531
rect 1468 467 1474 519
rect 1526 467 1532 519
rect 1468 459 1532 467
rect 1468 455 1484 459
rect 1518 455 1532 459
rect 1468 403 1474 455
rect 1526 403 1532 455
rect 1468 391 1532 403
rect 1468 339 1474 391
rect 1526 339 1532 391
rect 1468 327 1532 339
rect 1468 275 1474 327
rect 1526 275 1532 327
rect 1468 263 1532 275
rect 1468 211 1474 263
rect 1526 211 1532 263
rect 1468 209 1484 211
rect 1518 209 1532 211
rect 1468 199 1532 209
rect 1468 147 1474 199
rect 1526 147 1532 199
rect 1468 137 1484 147
rect 1518 137 1532 147
rect 1468 114 1532 137
rect 1566 517 1630 548
rect 1566 465 1572 517
rect 1624 465 1630 517
rect 1566 453 1630 465
rect 1566 401 1572 453
rect 1624 401 1630 453
rect 1566 389 1630 401
rect 1566 337 1572 389
rect 1624 337 1630 389
rect 1566 325 1630 337
rect 1566 273 1572 325
rect 1624 273 1630 325
rect 1566 261 1630 273
rect 1566 209 1572 261
rect 1624 209 1630 261
rect 1566 197 1630 209
rect 1566 145 1572 197
rect 1624 145 1630 197
rect 1566 114 1630 145
rect 1660 531 1724 552
rect 1660 519 1676 531
rect 1710 519 1724 531
rect 1660 467 1666 519
rect 1718 467 1724 519
rect 1660 459 1724 467
rect 1660 455 1676 459
rect 1710 455 1724 459
rect 1660 403 1666 455
rect 1718 403 1724 455
rect 1660 391 1724 403
rect 1660 339 1666 391
rect 1718 339 1724 391
rect 1660 327 1724 339
rect 1660 275 1666 327
rect 1718 275 1724 327
rect 1660 263 1724 275
rect 1660 211 1666 263
rect 1718 211 1724 263
rect 1660 209 1676 211
rect 1710 209 1724 211
rect 1660 199 1724 209
rect 1660 147 1666 199
rect 1718 147 1724 199
rect 1660 137 1676 147
rect 1710 137 1724 147
rect 1660 114 1724 137
rect 1758 517 1822 548
rect 1758 465 1764 517
rect 1816 465 1822 517
rect 1758 453 1822 465
rect 1758 401 1764 453
rect 1816 401 1822 453
rect 1758 389 1822 401
rect 1758 337 1764 389
rect 1816 337 1822 389
rect 1758 325 1822 337
rect 1758 273 1764 325
rect 1816 273 1822 325
rect 1758 261 1822 273
rect 1758 209 1764 261
rect 1816 209 1822 261
rect 1758 197 1822 209
rect 1758 145 1764 197
rect 1816 145 1822 197
rect 1758 114 1822 145
rect 78 26 1676 74
rect 82 -308 1680 -260
rect 34 -380 98 -344
rect 34 -432 40 -380
rect 92 -432 98 -380
rect 34 -444 98 -432
rect 34 -496 40 -444
rect 92 -496 98 -444
rect 34 -532 98 -496
rect 130 -379 194 -344
rect 130 -431 136 -379
rect 188 -431 194 -379
rect 130 -443 194 -431
rect 130 -495 136 -443
rect 188 -495 194 -443
rect 130 -530 194 -495
rect 226 -380 290 -344
rect 226 -432 232 -380
rect 284 -432 290 -380
rect 226 -444 290 -432
rect 226 -496 232 -444
rect 284 -496 290 -444
rect 226 -532 290 -496
rect 322 -379 386 -344
rect 322 -431 328 -379
rect 380 -431 386 -379
rect 322 -443 386 -431
rect 322 -495 328 -443
rect 380 -495 386 -443
rect 322 -530 386 -495
rect 418 -380 482 -344
rect 418 -432 424 -380
rect 476 -432 482 -380
rect 418 -444 482 -432
rect 418 -496 424 -444
rect 476 -496 482 -444
rect 418 -532 482 -496
rect 514 -379 578 -344
rect 514 -431 520 -379
rect 572 -431 578 -379
rect 514 -443 578 -431
rect 514 -495 520 -443
rect 572 -495 578 -443
rect 514 -530 578 -495
rect 610 -380 674 -344
rect 610 -432 616 -380
rect 668 -432 674 -380
rect 610 -444 674 -432
rect 610 -496 616 -444
rect 668 -496 674 -444
rect 610 -532 674 -496
rect 706 -379 770 -344
rect 706 -431 712 -379
rect 764 -431 770 -379
rect 706 -443 770 -431
rect 706 -495 712 -443
rect 764 -495 770 -443
rect 706 -530 770 -495
rect 802 -380 866 -344
rect 802 -432 808 -380
rect 860 -432 866 -380
rect 802 -444 866 -432
rect 802 -496 808 -444
rect 860 -496 866 -444
rect 802 -532 866 -496
rect 898 -379 962 -344
rect 898 -431 904 -379
rect 956 -431 962 -379
rect 898 -443 962 -431
rect 898 -495 904 -443
rect 956 -495 962 -443
rect 898 -530 962 -495
rect 994 -380 1058 -344
rect 994 -432 1000 -380
rect 1052 -432 1058 -380
rect 994 -444 1058 -432
rect 994 -496 1000 -444
rect 1052 -496 1058 -444
rect 994 -532 1058 -496
rect 1090 -379 1154 -344
rect 1090 -431 1096 -379
rect 1148 -431 1154 -379
rect 1090 -443 1154 -431
rect 1090 -495 1096 -443
rect 1148 -495 1154 -443
rect 1090 -530 1154 -495
rect 1186 -380 1250 -344
rect 1186 -432 1192 -380
rect 1244 -432 1250 -380
rect 1186 -444 1250 -432
rect 1186 -496 1192 -444
rect 1244 -496 1250 -444
rect 1186 -532 1250 -496
rect 1282 -379 1346 -344
rect 1282 -431 1288 -379
rect 1340 -431 1346 -379
rect 1282 -443 1346 -431
rect 1282 -495 1288 -443
rect 1340 -495 1346 -443
rect 1282 -530 1346 -495
rect 1378 -380 1442 -344
rect 1378 -432 1384 -380
rect 1436 -432 1442 -380
rect 1378 -444 1442 -432
rect 1378 -496 1384 -444
rect 1436 -496 1442 -444
rect 1378 -532 1442 -496
rect 1474 -379 1538 -344
rect 1474 -431 1480 -379
rect 1532 -431 1538 -379
rect 1474 -443 1538 -431
rect 1474 -495 1480 -443
rect 1532 -495 1538 -443
rect 1474 -530 1538 -495
rect 1570 -380 1634 -344
rect 1570 -432 1576 -380
rect 1628 -432 1634 -380
rect 1570 -444 1634 -432
rect 1570 -496 1576 -444
rect 1628 -496 1634 -444
rect 1570 -532 1634 -496
rect 1666 -379 1730 -344
rect 1666 -431 1672 -379
rect 1724 -431 1730 -379
rect 1666 -443 1730 -431
rect 1666 -495 1672 -443
rect 1724 -495 1730 -443
rect 1666 -530 1730 -495
rect 1762 -380 1826 -344
rect 1762 -432 1768 -380
rect 1820 -432 1826 -380
rect 1762 -444 1826 -432
rect 1762 -496 1768 -444
rect 1820 -496 1826 -444
rect 1762 -532 1826 -496
rect -166 -714 1776 -564
rect -163 -718 1776 -714
rect 34 -788 98 -752
rect 34 -840 40 -788
rect 92 -840 98 -788
rect 34 -852 98 -840
rect 34 -904 40 -852
rect 92 -904 98 -852
rect 34 -940 98 -904
rect 130 -789 194 -754
rect 130 -841 136 -789
rect 188 -841 194 -789
rect 130 -853 194 -841
rect 130 -905 136 -853
rect 188 -905 194 -853
rect 130 -940 194 -905
rect 226 -788 290 -752
rect 226 -840 232 -788
rect 284 -840 290 -788
rect 226 -852 290 -840
rect 226 -904 232 -852
rect 284 -904 290 -852
rect 226 -940 290 -904
rect 322 -789 386 -754
rect 322 -841 328 -789
rect 380 -841 386 -789
rect 322 -853 386 -841
rect 322 -905 328 -853
rect 380 -905 386 -853
rect 322 -940 386 -905
rect 418 -788 482 -752
rect 418 -840 424 -788
rect 476 -840 482 -788
rect 418 -852 482 -840
rect 418 -904 424 -852
rect 476 -904 482 -852
rect 418 -940 482 -904
rect 514 -789 578 -754
rect 514 -841 520 -789
rect 572 -841 578 -789
rect 514 -853 578 -841
rect 514 -905 520 -853
rect 572 -905 578 -853
rect 514 -940 578 -905
rect 610 -788 674 -752
rect 610 -840 616 -788
rect 668 -840 674 -788
rect 610 -852 674 -840
rect 610 -904 616 -852
rect 668 -904 674 -852
rect 610 -940 674 -904
rect 706 -789 770 -754
rect 706 -841 712 -789
rect 764 -841 770 -789
rect 706 -853 770 -841
rect 706 -905 712 -853
rect 764 -905 770 -853
rect 706 -940 770 -905
rect 802 -788 866 -752
rect 802 -840 808 -788
rect 860 -840 866 -788
rect 802 -852 866 -840
rect 802 -904 808 -852
rect 860 -904 866 -852
rect 802 -940 866 -904
rect 898 -789 962 -754
rect 898 -841 904 -789
rect 956 -841 962 -789
rect 898 -853 962 -841
rect 898 -905 904 -853
rect 956 -905 962 -853
rect 898 -940 962 -905
rect 994 -788 1058 -752
rect 994 -840 1000 -788
rect 1052 -840 1058 -788
rect 994 -852 1058 -840
rect 994 -904 1000 -852
rect 1052 -904 1058 -852
rect 994 -940 1058 -904
rect 1090 -789 1154 -754
rect 1090 -841 1096 -789
rect 1148 -841 1154 -789
rect 1090 -853 1154 -841
rect 1090 -905 1096 -853
rect 1148 -905 1154 -853
rect 1090 -940 1154 -905
rect 1186 -788 1250 -752
rect 1186 -840 1192 -788
rect 1244 -840 1250 -788
rect 1186 -852 1250 -840
rect 1186 -904 1192 -852
rect 1244 -904 1250 -852
rect 1186 -940 1250 -904
rect 1282 -789 1346 -754
rect 1282 -841 1288 -789
rect 1340 -841 1346 -789
rect 1282 -853 1346 -841
rect 1282 -905 1288 -853
rect 1340 -905 1346 -853
rect 1282 -940 1346 -905
rect 1378 -788 1442 -752
rect 1378 -840 1384 -788
rect 1436 -840 1442 -788
rect 1378 -852 1442 -840
rect 1378 -904 1384 -852
rect 1436 -904 1442 -852
rect 1378 -940 1442 -904
rect 1474 -789 1538 -754
rect 1474 -841 1480 -789
rect 1532 -841 1538 -789
rect 1474 -853 1538 -841
rect 1474 -905 1480 -853
rect 1532 -905 1538 -853
rect 1474 -940 1538 -905
rect 1570 -788 1634 -752
rect 1570 -840 1576 -788
rect 1628 -840 1634 -788
rect 1570 -852 1634 -840
rect 1570 -904 1576 -852
rect 1628 -904 1634 -852
rect 1570 -940 1634 -904
rect 1666 -789 1730 -754
rect 1666 -841 1672 -789
rect 1724 -841 1730 -789
rect 1666 -853 1730 -841
rect 1666 -905 1672 -853
rect 1724 -905 1730 -853
rect 1666 -940 1730 -905
rect 1762 -788 1826 -752
rect 1762 -840 1768 -788
rect 1820 -840 1826 -788
rect 1762 -852 1826 -840
rect 1762 -904 1768 -852
rect 1820 -904 1826 -852
rect 1762 -940 1826 -904
rect 80 -1022 1730 -974
rect -76 -1148 1924 -1142
rect -76 -1168 1926 -1148
rect -76 -1220 -57 -1168
rect -5 -1181 7 -1168
rect 59 -1181 71 -1168
rect 123 -1181 135 -1168
rect 187 -1181 199 -1168
rect 187 -1215 191 -1181
rect -5 -1220 7 -1215
rect 59 -1220 71 -1215
rect 123 -1220 135 -1215
rect 187 -1220 199 -1215
rect 251 -1220 263 -1168
rect 315 -1220 327 -1168
rect 379 -1220 391 -1168
rect 443 -1220 455 -1168
rect 507 -1181 519 -1168
rect 571 -1181 583 -1168
rect 635 -1181 647 -1168
rect 699 -1181 711 -1168
rect 763 -1181 775 -1168
rect 513 -1215 519 -1181
rect 763 -1215 767 -1181
rect 507 -1220 519 -1215
rect 571 -1220 583 -1215
rect 635 -1220 647 -1215
rect 699 -1220 711 -1215
rect 763 -1220 775 -1215
rect 827 -1220 839 -1168
rect 891 -1220 903 -1168
rect 955 -1220 967 -1168
rect 1019 -1220 1031 -1168
rect 1083 -1181 1095 -1168
rect 1147 -1181 1159 -1168
rect 1211 -1181 1223 -1168
rect 1275 -1181 1287 -1168
rect 1339 -1181 1351 -1168
rect 1089 -1215 1095 -1181
rect 1339 -1215 1343 -1181
rect 1083 -1220 1095 -1215
rect 1147 -1220 1159 -1215
rect 1211 -1220 1223 -1215
rect 1275 -1220 1287 -1215
rect 1339 -1220 1351 -1215
rect 1403 -1220 1415 -1168
rect 1467 -1220 1479 -1168
rect 1531 -1220 1543 -1168
rect 1595 -1220 1607 -1168
rect 1659 -1181 1671 -1168
rect 1723 -1181 1735 -1168
rect 1787 -1181 1799 -1168
rect 1851 -1181 1863 -1168
rect 1665 -1215 1671 -1181
rect 1659 -1220 1671 -1215
rect 1723 -1220 1735 -1215
rect 1787 -1220 1799 -1215
rect 1851 -1220 1863 -1215
rect 1915 -1220 1926 -1168
rect -76 -1234 1926 -1220
rect -74 -1246 1926 -1234
<< via1 >>
rect -66 1522 -14 1536
rect -66 1488 -33 1522
rect -33 1488 -14 1522
rect -66 1484 -14 1488
rect -2 1522 50 1536
rect -2 1488 5 1522
rect 5 1488 39 1522
rect 39 1488 50 1522
rect -2 1484 50 1488
rect 62 1522 114 1536
rect 62 1488 77 1522
rect 77 1488 111 1522
rect 111 1488 114 1522
rect 62 1484 114 1488
rect 126 1522 178 1536
rect 190 1522 242 1536
rect 254 1522 306 1536
rect 318 1522 370 1536
rect 382 1522 434 1536
rect 446 1522 498 1536
rect 510 1522 562 1536
rect 126 1488 149 1522
rect 149 1488 178 1522
rect 190 1488 221 1522
rect 221 1488 242 1522
rect 254 1488 255 1522
rect 255 1488 293 1522
rect 293 1488 306 1522
rect 318 1488 327 1522
rect 327 1488 365 1522
rect 365 1488 370 1522
rect 382 1488 399 1522
rect 399 1488 434 1522
rect 446 1488 471 1522
rect 471 1488 498 1522
rect 510 1488 543 1522
rect 543 1488 562 1522
rect 126 1484 178 1488
rect 190 1484 242 1488
rect 254 1484 306 1488
rect 318 1484 370 1488
rect 382 1484 434 1488
rect 446 1484 498 1488
rect 510 1484 562 1488
rect 574 1522 626 1536
rect 574 1488 581 1522
rect 581 1488 615 1522
rect 615 1488 626 1522
rect 574 1484 626 1488
rect 638 1522 690 1536
rect 638 1488 653 1522
rect 653 1488 687 1522
rect 687 1488 690 1522
rect 638 1484 690 1488
rect 702 1522 754 1536
rect 766 1522 818 1536
rect 830 1522 882 1536
rect 894 1522 946 1536
rect 958 1522 1010 1536
rect 1022 1522 1074 1536
rect 1086 1522 1138 1536
rect 702 1488 725 1522
rect 725 1488 754 1522
rect 766 1488 797 1522
rect 797 1488 818 1522
rect 830 1488 831 1522
rect 831 1488 869 1522
rect 869 1488 882 1522
rect 894 1488 903 1522
rect 903 1488 941 1522
rect 941 1488 946 1522
rect 958 1488 975 1522
rect 975 1488 1010 1522
rect 1022 1488 1047 1522
rect 1047 1488 1074 1522
rect 1086 1488 1119 1522
rect 1119 1488 1138 1522
rect 702 1484 754 1488
rect 766 1484 818 1488
rect 830 1484 882 1488
rect 894 1484 946 1488
rect 958 1484 1010 1488
rect 1022 1484 1074 1488
rect 1086 1484 1138 1488
rect 1150 1522 1202 1536
rect 1150 1488 1157 1522
rect 1157 1488 1191 1522
rect 1191 1488 1202 1522
rect 1150 1484 1202 1488
rect 1214 1522 1266 1536
rect 1214 1488 1229 1522
rect 1229 1488 1263 1522
rect 1263 1488 1266 1522
rect 1214 1484 1266 1488
rect 1278 1522 1330 1536
rect 1342 1522 1394 1536
rect 1406 1522 1458 1536
rect 1470 1522 1522 1536
rect 1534 1522 1586 1536
rect 1598 1522 1650 1536
rect 1662 1522 1714 1536
rect 1278 1488 1301 1522
rect 1301 1488 1330 1522
rect 1342 1488 1373 1522
rect 1373 1488 1394 1522
rect 1406 1488 1407 1522
rect 1407 1488 1445 1522
rect 1445 1488 1458 1522
rect 1470 1488 1479 1522
rect 1479 1488 1517 1522
rect 1517 1488 1522 1522
rect 1534 1488 1551 1522
rect 1551 1488 1586 1522
rect 1598 1488 1623 1522
rect 1623 1488 1650 1522
rect 1662 1488 1695 1522
rect 1695 1488 1714 1522
rect 1278 1484 1330 1488
rect 1342 1484 1394 1488
rect 1406 1484 1458 1488
rect 1470 1484 1522 1488
rect 1534 1484 1586 1488
rect 1598 1484 1650 1488
rect 1662 1484 1714 1488
rect 1726 1522 1778 1536
rect 1726 1488 1733 1522
rect 1733 1488 1767 1522
rect 1767 1488 1778 1522
rect 1726 1484 1778 1488
rect 1790 1522 1842 1536
rect 1790 1488 1805 1522
rect 1805 1488 1839 1522
rect 1839 1488 1842 1522
rect 1790 1484 1842 1488
rect 1854 1522 1906 1536
rect 1854 1488 1877 1522
rect 1877 1488 1906 1522
rect 1854 1484 1906 1488
rect 36 1143 88 1195
rect 36 1079 88 1131
rect 36 1015 88 1067
rect 36 951 88 1003
rect 36 887 88 939
rect 36 823 88 875
rect 130 1175 140 1197
rect 140 1175 174 1197
rect 174 1175 182 1197
rect 130 1145 182 1175
rect 130 1103 140 1133
rect 140 1103 174 1133
rect 174 1103 182 1133
rect 130 1081 182 1103
rect 130 1065 182 1069
rect 130 1031 140 1065
rect 140 1031 174 1065
rect 174 1031 182 1065
rect 130 1017 182 1031
rect 130 993 182 1005
rect 130 959 140 993
rect 140 959 174 993
rect 174 959 182 993
rect 130 953 182 959
rect 130 921 182 941
rect 130 889 140 921
rect 140 889 174 921
rect 174 889 182 921
rect 130 849 182 877
rect 130 825 140 849
rect 140 825 174 849
rect 174 825 182 849
rect 228 1143 280 1195
rect 228 1079 280 1131
rect 228 1015 280 1067
rect 228 951 280 1003
rect 228 887 280 939
rect 228 823 280 875
rect 322 1175 332 1197
rect 332 1175 366 1197
rect 366 1175 374 1197
rect 322 1145 374 1175
rect 322 1103 332 1133
rect 332 1103 366 1133
rect 366 1103 374 1133
rect 322 1081 374 1103
rect 322 1065 374 1069
rect 322 1031 332 1065
rect 332 1031 366 1065
rect 366 1031 374 1065
rect 322 1017 374 1031
rect 322 993 374 1005
rect 322 959 332 993
rect 332 959 366 993
rect 366 959 374 993
rect 322 953 374 959
rect 322 921 374 941
rect 322 889 332 921
rect 332 889 366 921
rect 366 889 374 921
rect 322 849 374 877
rect 322 825 332 849
rect 332 825 366 849
rect 366 825 374 849
rect 420 1143 472 1195
rect 420 1079 472 1131
rect 420 1015 472 1067
rect 420 951 472 1003
rect 420 887 472 939
rect 420 823 472 875
rect 514 1175 524 1197
rect 524 1175 558 1197
rect 558 1175 566 1197
rect 514 1145 566 1175
rect 514 1103 524 1133
rect 524 1103 558 1133
rect 558 1103 566 1133
rect 514 1081 566 1103
rect 514 1065 566 1069
rect 514 1031 524 1065
rect 524 1031 558 1065
rect 558 1031 566 1065
rect 514 1017 566 1031
rect 514 993 566 1005
rect 514 959 524 993
rect 524 959 558 993
rect 558 959 566 993
rect 514 953 566 959
rect 514 921 566 941
rect 514 889 524 921
rect 524 889 558 921
rect 558 889 566 921
rect 514 849 566 877
rect 514 825 524 849
rect 524 825 558 849
rect 558 825 566 849
rect 612 1143 664 1195
rect 612 1079 664 1131
rect 612 1015 664 1067
rect 612 951 664 1003
rect 612 887 664 939
rect 612 823 664 875
rect 706 1175 716 1197
rect 716 1175 750 1197
rect 750 1175 758 1197
rect 706 1145 758 1175
rect 706 1103 716 1133
rect 716 1103 750 1133
rect 750 1103 758 1133
rect 706 1081 758 1103
rect 706 1065 758 1069
rect 706 1031 716 1065
rect 716 1031 750 1065
rect 750 1031 758 1065
rect 706 1017 758 1031
rect 706 993 758 1005
rect 706 959 716 993
rect 716 959 750 993
rect 750 959 758 993
rect 706 953 758 959
rect 706 921 758 941
rect 706 889 716 921
rect 716 889 750 921
rect 750 889 758 921
rect 706 849 758 877
rect 706 825 716 849
rect 716 825 750 849
rect 750 825 758 849
rect 804 1143 856 1195
rect 804 1079 856 1131
rect 804 1015 856 1067
rect 804 951 856 1003
rect 804 887 856 939
rect 804 823 856 875
rect 898 1175 908 1197
rect 908 1175 942 1197
rect 942 1175 950 1197
rect 898 1145 950 1175
rect 898 1103 908 1133
rect 908 1103 942 1133
rect 942 1103 950 1133
rect 898 1081 950 1103
rect 898 1065 950 1069
rect 898 1031 908 1065
rect 908 1031 942 1065
rect 942 1031 950 1065
rect 898 1017 950 1031
rect 898 993 950 1005
rect 898 959 908 993
rect 908 959 942 993
rect 942 959 950 993
rect 898 953 950 959
rect 898 921 950 941
rect 898 889 908 921
rect 908 889 942 921
rect 942 889 950 921
rect 898 849 950 877
rect 898 825 908 849
rect 908 825 942 849
rect 942 825 950 849
rect 996 1143 1048 1195
rect 996 1079 1048 1131
rect 996 1015 1048 1067
rect 996 951 1048 1003
rect 996 887 1048 939
rect 996 823 1048 875
rect 1090 1175 1100 1197
rect 1100 1175 1134 1197
rect 1134 1175 1142 1197
rect 1090 1145 1142 1175
rect 1090 1103 1100 1133
rect 1100 1103 1134 1133
rect 1134 1103 1142 1133
rect 1090 1081 1142 1103
rect 1090 1065 1142 1069
rect 1090 1031 1100 1065
rect 1100 1031 1134 1065
rect 1134 1031 1142 1065
rect 1090 1017 1142 1031
rect 1090 993 1142 1005
rect 1090 959 1100 993
rect 1100 959 1134 993
rect 1134 959 1142 993
rect 1090 953 1142 959
rect 1090 921 1142 941
rect 1090 889 1100 921
rect 1100 889 1134 921
rect 1134 889 1142 921
rect 1090 849 1142 877
rect 1090 825 1100 849
rect 1100 825 1134 849
rect 1134 825 1142 849
rect 1188 1143 1240 1195
rect 1188 1079 1240 1131
rect 1188 1015 1240 1067
rect 1188 951 1240 1003
rect 1188 887 1240 939
rect 1188 823 1240 875
rect 1282 1175 1292 1197
rect 1292 1175 1326 1197
rect 1326 1175 1334 1197
rect 1282 1145 1334 1175
rect 1282 1103 1292 1133
rect 1292 1103 1326 1133
rect 1326 1103 1334 1133
rect 1282 1081 1334 1103
rect 1282 1065 1334 1069
rect 1282 1031 1292 1065
rect 1292 1031 1326 1065
rect 1326 1031 1334 1065
rect 1282 1017 1334 1031
rect 1282 993 1334 1005
rect 1282 959 1292 993
rect 1292 959 1326 993
rect 1326 959 1334 993
rect 1282 953 1334 959
rect 1282 921 1334 941
rect 1282 889 1292 921
rect 1292 889 1326 921
rect 1326 889 1334 921
rect 1282 849 1334 877
rect 1282 825 1292 849
rect 1292 825 1326 849
rect 1326 825 1334 849
rect 1380 1143 1432 1195
rect 1380 1079 1432 1131
rect 1380 1015 1432 1067
rect 1380 951 1432 1003
rect 1380 887 1432 939
rect 1380 823 1432 875
rect 1474 1175 1484 1197
rect 1484 1175 1518 1197
rect 1518 1175 1526 1197
rect 1474 1145 1526 1175
rect 1474 1103 1484 1133
rect 1484 1103 1518 1133
rect 1518 1103 1526 1133
rect 1474 1081 1526 1103
rect 1474 1065 1526 1069
rect 1474 1031 1484 1065
rect 1484 1031 1518 1065
rect 1518 1031 1526 1065
rect 1474 1017 1526 1031
rect 1474 993 1526 1005
rect 1474 959 1484 993
rect 1484 959 1518 993
rect 1518 959 1526 993
rect 1474 953 1526 959
rect 1474 921 1526 941
rect 1474 889 1484 921
rect 1484 889 1518 921
rect 1518 889 1526 921
rect 1474 849 1526 877
rect 1474 825 1484 849
rect 1484 825 1518 849
rect 1518 825 1526 849
rect 1572 1143 1624 1195
rect 1572 1079 1624 1131
rect 1572 1015 1624 1067
rect 1572 951 1624 1003
rect 1572 887 1624 939
rect 1572 823 1624 875
rect 1666 1175 1676 1197
rect 1676 1175 1710 1197
rect 1710 1175 1718 1197
rect 1666 1145 1718 1175
rect 1666 1103 1676 1133
rect 1676 1103 1710 1133
rect 1710 1103 1718 1133
rect 1666 1081 1718 1103
rect 1666 1065 1718 1069
rect 1666 1031 1676 1065
rect 1676 1031 1710 1065
rect 1710 1031 1718 1065
rect 1666 1017 1718 1031
rect 1666 993 1718 1005
rect 1666 959 1676 993
rect 1676 959 1710 993
rect 1710 959 1718 993
rect 1666 953 1718 959
rect 1666 921 1718 941
rect 1666 889 1676 921
rect 1676 889 1710 921
rect 1710 889 1718 921
rect 1666 849 1718 877
rect 1666 825 1676 849
rect 1676 825 1710 849
rect 1710 825 1718 849
rect 1764 1143 1816 1195
rect 1764 1079 1816 1131
rect 1764 1015 1816 1067
rect 1764 951 1816 1003
rect 1764 887 1816 939
rect 1764 823 1816 875
rect 36 465 88 517
rect 36 401 88 453
rect 36 337 88 389
rect 36 273 88 325
rect 36 209 88 261
rect 36 145 88 197
rect 130 497 140 519
rect 140 497 174 519
rect 174 497 182 519
rect 130 467 182 497
rect 130 425 140 455
rect 140 425 174 455
rect 174 425 182 455
rect 130 403 182 425
rect 130 387 182 391
rect 130 353 140 387
rect 140 353 174 387
rect 174 353 182 387
rect 130 339 182 353
rect 130 315 182 327
rect 130 281 140 315
rect 140 281 174 315
rect 174 281 182 315
rect 130 275 182 281
rect 130 243 182 263
rect 130 211 140 243
rect 140 211 174 243
rect 174 211 182 243
rect 130 171 182 199
rect 130 147 140 171
rect 140 147 174 171
rect 174 147 182 171
rect 228 465 280 517
rect 228 401 280 453
rect 228 337 280 389
rect 228 273 280 325
rect 228 209 280 261
rect 228 145 280 197
rect 322 497 332 519
rect 332 497 366 519
rect 366 497 374 519
rect 322 467 374 497
rect 322 425 332 455
rect 332 425 366 455
rect 366 425 374 455
rect 322 403 374 425
rect 322 387 374 391
rect 322 353 332 387
rect 332 353 366 387
rect 366 353 374 387
rect 322 339 374 353
rect 322 315 374 327
rect 322 281 332 315
rect 332 281 366 315
rect 366 281 374 315
rect 322 275 374 281
rect 322 243 374 263
rect 322 211 332 243
rect 332 211 366 243
rect 366 211 374 243
rect 322 171 374 199
rect 322 147 332 171
rect 332 147 366 171
rect 366 147 374 171
rect 420 465 472 517
rect 420 401 472 453
rect 420 337 472 389
rect 420 273 472 325
rect 420 209 472 261
rect 420 145 472 197
rect 514 497 524 519
rect 524 497 558 519
rect 558 497 566 519
rect 514 467 566 497
rect 514 425 524 455
rect 524 425 558 455
rect 558 425 566 455
rect 514 403 566 425
rect 514 387 566 391
rect 514 353 524 387
rect 524 353 558 387
rect 558 353 566 387
rect 514 339 566 353
rect 514 315 566 327
rect 514 281 524 315
rect 524 281 558 315
rect 558 281 566 315
rect 514 275 566 281
rect 514 243 566 263
rect 514 211 524 243
rect 524 211 558 243
rect 558 211 566 243
rect 514 171 566 199
rect 514 147 524 171
rect 524 147 558 171
rect 558 147 566 171
rect 612 465 664 517
rect 612 401 664 453
rect 612 337 664 389
rect 612 273 664 325
rect 612 209 664 261
rect 612 145 664 197
rect 706 497 716 519
rect 716 497 750 519
rect 750 497 758 519
rect 706 467 758 497
rect 706 425 716 455
rect 716 425 750 455
rect 750 425 758 455
rect 706 403 758 425
rect 706 387 758 391
rect 706 353 716 387
rect 716 353 750 387
rect 750 353 758 387
rect 706 339 758 353
rect 706 315 758 327
rect 706 281 716 315
rect 716 281 750 315
rect 750 281 758 315
rect 706 275 758 281
rect 706 243 758 263
rect 706 211 716 243
rect 716 211 750 243
rect 750 211 758 243
rect 706 171 758 199
rect 706 147 716 171
rect 716 147 750 171
rect 750 147 758 171
rect 804 465 856 517
rect 804 401 856 453
rect 804 337 856 389
rect 804 273 856 325
rect 804 209 856 261
rect 804 145 856 197
rect 898 497 908 519
rect 908 497 942 519
rect 942 497 950 519
rect 898 467 950 497
rect 898 425 908 455
rect 908 425 942 455
rect 942 425 950 455
rect 898 403 950 425
rect 898 387 950 391
rect 898 353 908 387
rect 908 353 942 387
rect 942 353 950 387
rect 898 339 950 353
rect 898 315 950 327
rect 898 281 908 315
rect 908 281 942 315
rect 942 281 950 315
rect 898 275 950 281
rect 898 243 950 263
rect 898 211 908 243
rect 908 211 942 243
rect 942 211 950 243
rect 898 171 950 199
rect 898 147 908 171
rect 908 147 942 171
rect 942 147 950 171
rect 996 465 1048 517
rect 996 401 1048 453
rect 996 337 1048 389
rect 996 273 1048 325
rect 996 209 1048 261
rect 996 145 1048 197
rect 1090 497 1100 519
rect 1100 497 1134 519
rect 1134 497 1142 519
rect 1090 467 1142 497
rect 1090 425 1100 455
rect 1100 425 1134 455
rect 1134 425 1142 455
rect 1090 403 1142 425
rect 1090 387 1142 391
rect 1090 353 1100 387
rect 1100 353 1134 387
rect 1134 353 1142 387
rect 1090 339 1142 353
rect 1090 315 1142 327
rect 1090 281 1100 315
rect 1100 281 1134 315
rect 1134 281 1142 315
rect 1090 275 1142 281
rect 1090 243 1142 263
rect 1090 211 1100 243
rect 1100 211 1134 243
rect 1134 211 1142 243
rect 1090 171 1142 199
rect 1090 147 1100 171
rect 1100 147 1134 171
rect 1134 147 1142 171
rect 1188 465 1240 517
rect 1188 401 1240 453
rect 1188 337 1240 389
rect 1188 273 1240 325
rect 1188 209 1240 261
rect 1188 145 1240 197
rect 1282 497 1292 519
rect 1292 497 1326 519
rect 1326 497 1334 519
rect 1282 467 1334 497
rect 1282 425 1292 455
rect 1292 425 1326 455
rect 1326 425 1334 455
rect 1282 403 1334 425
rect 1282 387 1334 391
rect 1282 353 1292 387
rect 1292 353 1326 387
rect 1326 353 1334 387
rect 1282 339 1334 353
rect 1282 315 1334 327
rect 1282 281 1292 315
rect 1292 281 1326 315
rect 1326 281 1334 315
rect 1282 275 1334 281
rect 1282 243 1334 263
rect 1282 211 1292 243
rect 1292 211 1326 243
rect 1326 211 1334 243
rect 1282 171 1334 199
rect 1282 147 1292 171
rect 1292 147 1326 171
rect 1326 147 1334 171
rect 1380 465 1432 517
rect 1380 401 1432 453
rect 1380 337 1432 389
rect 1380 273 1432 325
rect 1380 209 1432 261
rect 1380 145 1432 197
rect 1474 497 1484 519
rect 1484 497 1518 519
rect 1518 497 1526 519
rect 1474 467 1526 497
rect 1474 425 1484 455
rect 1484 425 1518 455
rect 1518 425 1526 455
rect 1474 403 1526 425
rect 1474 387 1526 391
rect 1474 353 1484 387
rect 1484 353 1518 387
rect 1518 353 1526 387
rect 1474 339 1526 353
rect 1474 315 1526 327
rect 1474 281 1484 315
rect 1484 281 1518 315
rect 1518 281 1526 315
rect 1474 275 1526 281
rect 1474 243 1526 263
rect 1474 211 1484 243
rect 1484 211 1518 243
rect 1518 211 1526 243
rect 1474 171 1526 199
rect 1474 147 1484 171
rect 1484 147 1518 171
rect 1518 147 1526 171
rect 1572 465 1624 517
rect 1572 401 1624 453
rect 1572 337 1624 389
rect 1572 273 1624 325
rect 1572 209 1624 261
rect 1572 145 1624 197
rect 1666 497 1676 519
rect 1676 497 1710 519
rect 1710 497 1718 519
rect 1666 467 1718 497
rect 1666 425 1676 455
rect 1676 425 1710 455
rect 1710 425 1718 455
rect 1666 403 1718 425
rect 1666 387 1718 391
rect 1666 353 1676 387
rect 1676 353 1710 387
rect 1710 353 1718 387
rect 1666 339 1718 353
rect 1666 315 1718 327
rect 1666 281 1676 315
rect 1676 281 1710 315
rect 1710 281 1718 315
rect 1666 275 1718 281
rect 1666 243 1718 263
rect 1666 211 1676 243
rect 1676 211 1710 243
rect 1710 211 1718 243
rect 1666 171 1718 199
rect 1666 147 1676 171
rect 1676 147 1710 171
rect 1710 147 1718 171
rect 1764 465 1816 517
rect 1764 401 1816 453
rect 1764 337 1816 389
rect 1764 273 1816 325
rect 1764 209 1816 261
rect 1764 145 1816 197
rect 40 -432 92 -380
rect 40 -496 92 -444
rect 136 -431 188 -379
rect 136 -495 188 -443
rect 232 -432 284 -380
rect 232 -496 284 -444
rect 328 -431 380 -379
rect 328 -495 380 -443
rect 424 -432 476 -380
rect 424 -496 476 -444
rect 520 -431 572 -379
rect 520 -495 572 -443
rect 616 -432 668 -380
rect 616 -496 668 -444
rect 712 -431 764 -379
rect 712 -495 764 -443
rect 808 -432 860 -380
rect 808 -496 860 -444
rect 904 -431 956 -379
rect 904 -495 956 -443
rect 1000 -432 1052 -380
rect 1000 -496 1052 -444
rect 1096 -431 1148 -379
rect 1096 -495 1148 -443
rect 1192 -432 1244 -380
rect 1192 -496 1244 -444
rect 1288 -431 1340 -379
rect 1288 -495 1340 -443
rect 1384 -432 1436 -380
rect 1384 -496 1436 -444
rect 1480 -431 1532 -379
rect 1480 -495 1532 -443
rect 1576 -432 1628 -380
rect 1576 -496 1628 -444
rect 1672 -431 1724 -379
rect 1672 -495 1724 -443
rect 1768 -432 1820 -380
rect 1768 -496 1820 -444
rect 40 -840 92 -788
rect 40 -904 92 -852
rect 136 -841 188 -789
rect 136 -905 188 -853
rect 232 -840 284 -788
rect 232 -904 284 -852
rect 328 -841 380 -789
rect 328 -905 380 -853
rect 424 -840 476 -788
rect 424 -904 476 -852
rect 520 -841 572 -789
rect 520 -905 572 -853
rect 616 -840 668 -788
rect 616 -904 668 -852
rect 712 -841 764 -789
rect 712 -905 764 -853
rect 808 -840 860 -788
rect 808 -904 860 -852
rect 904 -841 956 -789
rect 904 -905 956 -853
rect 1000 -840 1052 -788
rect 1000 -904 1052 -852
rect 1096 -841 1148 -789
rect 1096 -905 1148 -853
rect 1192 -840 1244 -788
rect 1192 -904 1244 -852
rect 1288 -841 1340 -789
rect 1288 -905 1340 -853
rect 1384 -840 1436 -788
rect 1384 -904 1436 -852
rect 1480 -841 1532 -789
rect 1480 -905 1532 -853
rect 1576 -840 1628 -788
rect 1576 -904 1628 -852
rect 1672 -841 1724 -789
rect 1672 -905 1724 -853
rect 1768 -840 1820 -788
rect 1768 -904 1820 -852
rect -57 -1181 -5 -1168
rect 7 -1181 59 -1168
rect 71 -1181 123 -1168
rect 135 -1181 187 -1168
rect 199 -1181 251 -1168
rect -57 -1215 -25 -1181
rect -25 -1215 -5 -1181
rect 7 -1215 9 -1181
rect 9 -1215 47 -1181
rect 47 -1215 59 -1181
rect 71 -1215 81 -1181
rect 81 -1215 119 -1181
rect 119 -1215 123 -1181
rect 135 -1215 153 -1181
rect 153 -1215 187 -1181
rect 199 -1215 225 -1181
rect 225 -1215 251 -1181
rect -57 -1220 -5 -1215
rect 7 -1220 59 -1215
rect 71 -1220 123 -1215
rect 135 -1220 187 -1215
rect 199 -1220 251 -1215
rect 263 -1181 315 -1168
rect 263 -1215 297 -1181
rect 297 -1215 315 -1181
rect 263 -1220 315 -1215
rect 327 -1181 379 -1168
rect 327 -1215 335 -1181
rect 335 -1215 369 -1181
rect 369 -1215 379 -1181
rect 327 -1220 379 -1215
rect 391 -1181 443 -1168
rect 391 -1215 407 -1181
rect 407 -1215 441 -1181
rect 441 -1215 443 -1181
rect 391 -1220 443 -1215
rect 455 -1181 507 -1168
rect 519 -1181 571 -1168
rect 583 -1181 635 -1168
rect 647 -1181 699 -1168
rect 711 -1181 763 -1168
rect 775 -1181 827 -1168
rect 455 -1215 479 -1181
rect 479 -1215 507 -1181
rect 519 -1215 551 -1181
rect 551 -1215 571 -1181
rect 583 -1215 585 -1181
rect 585 -1215 623 -1181
rect 623 -1215 635 -1181
rect 647 -1215 657 -1181
rect 657 -1215 695 -1181
rect 695 -1215 699 -1181
rect 711 -1215 729 -1181
rect 729 -1215 763 -1181
rect 775 -1215 801 -1181
rect 801 -1215 827 -1181
rect 455 -1220 507 -1215
rect 519 -1220 571 -1215
rect 583 -1220 635 -1215
rect 647 -1220 699 -1215
rect 711 -1220 763 -1215
rect 775 -1220 827 -1215
rect 839 -1181 891 -1168
rect 839 -1215 873 -1181
rect 873 -1215 891 -1181
rect 839 -1220 891 -1215
rect 903 -1181 955 -1168
rect 903 -1215 911 -1181
rect 911 -1215 945 -1181
rect 945 -1215 955 -1181
rect 903 -1220 955 -1215
rect 967 -1181 1019 -1168
rect 967 -1215 983 -1181
rect 983 -1215 1017 -1181
rect 1017 -1215 1019 -1181
rect 967 -1220 1019 -1215
rect 1031 -1181 1083 -1168
rect 1095 -1181 1147 -1168
rect 1159 -1181 1211 -1168
rect 1223 -1181 1275 -1168
rect 1287 -1181 1339 -1168
rect 1351 -1181 1403 -1168
rect 1031 -1215 1055 -1181
rect 1055 -1215 1083 -1181
rect 1095 -1215 1127 -1181
rect 1127 -1215 1147 -1181
rect 1159 -1215 1161 -1181
rect 1161 -1215 1199 -1181
rect 1199 -1215 1211 -1181
rect 1223 -1215 1233 -1181
rect 1233 -1215 1271 -1181
rect 1271 -1215 1275 -1181
rect 1287 -1215 1305 -1181
rect 1305 -1215 1339 -1181
rect 1351 -1215 1377 -1181
rect 1377 -1215 1403 -1181
rect 1031 -1220 1083 -1215
rect 1095 -1220 1147 -1215
rect 1159 -1220 1211 -1215
rect 1223 -1220 1275 -1215
rect 1287 -1220 1339 -1215
rect 1351 -1220 1403 -1215
rect 1415 -1181 1467 -1168
rect 1415 -1215 1449 -1181
rect 1449 -1215 1467 -1181
rect 1415 -1220 1467 -1215
rect 1479 -1181 1531 -1168
rect 1479 -1215 1487 -1181
rect 1487 -1215 1521 -1181
rect 1521 -1215 1531 -1181
rect 1479 -1220 1531 -1215
rect 1543 -1181 1595 -1168
rect 1543 -1215 1559 -1181
rect 1559 -1215 1593 -1181
rect 1593 -1215 1595 -1181
rect 1543 -1220 1595 -1215
rect 1607 -1181 1659 -1168
rect 1671 -1181 1723 -1168
rect 1735 -1181 1787 -1168
rect 1799 -1181 1851 -1168
rect 1863 -1181 1915 -1168
rect 1607 -1215 1631 -1181
rect 1631 -1215 1659 -1181
rect 1671 -1215 1703 -1181
rect 1703 -1215 1723 -1181
rect 1735 -1215 1737 -1181
rect 1737 -1215 1775 -1181
rect 1775 -1215 1787 -1181
rect 1799 -1215 1809 -1181
rect 1809 -1215 1847 -1181
rect 1847 -1215 1851 -1181
rect 1863 -1215 1881 -1181
rect 1881 -1215 1915 -1181
rect 1607 -1220 1659 -1215
rect 1671 -1220 1723 -1215
rect 1735 -1220 1787 -1215
rect 1799 -1220 1851 -1215
rect 1863 -1220 1915 -1215
<< metal2 >>
rect -106 1536 1956 1598
rect -106 1484 -66 1536
rect -14 1484 -2 1536
rect 50 1484 62 1536
rect 114 1484 126 1536
rect 178 1484 190 1536
rect 242 1484 254 1536
rect 306 1484 318 1536
rect 370 1484 382 1536
rect 434 1484 446 1536
rect 498 1484 510 1536
rect 562 1484 574 1536
rect 626 1484 638 1536
rect 690 1484 702 1536
rect 754 1484 766 1536
rect 818 1484 830 1536
rect 882 1484 894 1536
rect 946 1484 958 1536
rect 1010 1484 1022 1536
rect 1074 1484 1086 1536
rect 1138 1484 1150 1536
rect 1202 1484 1214 1536
rect 1266 1484 1278 1536
rect 1330 1484 1342 1536
rect 1394 1484 1406 1536
rect 1458 1484 1470 1536
rect 1522 1484 1534 1536
rect 1586 1484 1598 1536
rect 1650 1484 1662 1536
rect 1714 1484 1726 1536
rect 1778 1484 1790 1536
rect 1842 1484 1854 1536
rect 1906 1484 1956 1536
rect -106 1470 1956 1484
rect 30 1196 94 1226
rect 30 1140 34 1196
rect 90 1140 94 1196
rect 30 1131 94 1140
rect 30 1116 36 1131
rect 88 1116 94 1131
rect 30 1060 34 1116
rect 90 1060 94 1116
rect 30 1036 36 1060
rect 88 1036 94 1060
rect 30 980 34 1036
rect 90 980 94 1036
rect 30 956 36 980
rect 88 956 94 980
rect 30 900 34 956
rect 90 900 94 956
rect 30 887 36 900
rect 88 887 94 900
rect 30 876 94 887
rect 30 820 34 876
rect 90 820 94 876
rect 30 792 94 820
rect 124 1197 188 1470
rect 124 1145 130 1197
rect 182 1145 188 1197
rect 124 1133 188 1145
rect 124 1081 130 1133
rect 182 1081 188 1133
rect 124 1069 188 1081
rect 124 1017 130 1069
rect 182 1017 188 1069
rect 124 1005 188 1017
rect 124 953 130 1005
rect 182 953 188 1005
rect 124 941 188 953
rect 124 889 130 941
rect 182 889 188 941
rect 124 877 188 889
rect 124 825 130 877
rect 182 825 188 877
rect 30 518 94 548
rect 30 462 34 518
rect 90 462 94 518
rect 30 453 94 462
rect 30 438 36 453
rect 88 438 94 453
rect 30 382 34 438
rect 90 382 94 438
rect 30 358 36 382
rect 88 358 94 382
rect 30 302 34 358
rect 90 302 94 358
rect 30 278 36 302
rect 88 278 94 302
rect 30 222 34 278
rect 90 222 94 278
rect 30 209 36 222
rect 88 209 94 222
rect 30 198 94 209
rect 30 142 34 198
rect 90 142 94 198
rect 30 114 94 142
rect 124 519 188 825
rect 222 1196 286 1226
rect 222 1140 226 1196
rect 282 1140 286 1196
rect 222 1131 286 1140
rect 222 1116 228 1131
rect 280 1116 286 1131
rect 222 1060 226 1116
rect 282 1060 286 1116
rect 222 1036 228 1060
rect 280 1036 286 1060
rect 222 980 226 1036
rect 282 980 286 1036
rect 222 956 228 980
rect 280 956 286 980
rect 222 900 226 956
rect 282 900 286 956
rect 222 887 228 900
rect 280 887 286 900
rect 222 876 286 887
rect 222 820 226 876
rect 282 820 286 876
rect 222 792 286 820
rect 316 1197 380 1470
rect 508 1462 1242 1470
rect 316 1145 322 1197
rect 374 1145 380 1197
rect 316 1133 380 1145
rect 316 1081 322 1133
rect 374 1081 380 1133
rect 316 1069 380 1081
rect 316 1017 322 1069
rect 374 1017 380 1069
rect 316 1005 380 1017
rect 316 953 322 1005
rect 374 953 380 1005
rect 316 941 380 953
rect 316 889 322 941
rect 374 889 380 941
rect 316 877 380 889
rect 316 825 322 877
rect 374 825 380 877
rect 124 467 130 519
rect 182 467 188 519
rect 124 455 188 467
rect 124 403 130 455
rect 182 403 188 455
rect 124 391 188 403
rect 124 339 130 391
rect 182 339 188 391
rect 124 327 188 339
rect 124 275 130 327
rect 182 275 188 327
rect 124 263 188 275
rect 124 211 130 263
rect 182 211 188 263
rect 124 199 188 211
rect 124 147 130 199
rect 182 147 188 199
rect 124 114 188 147
rect 222 518 286 548
rect 222 462 226 518
rect 282 462 286 518
rect 222 453 286 462
rect 222 438 228 453
rect 280 438 286 453
rect 222 382 226 438
rect 282 382 286 438
rect 222 358 228 382
rect 280 358 286 382
rect 222 302 226 358
rect 282 302 286 358
rect 222 278 228 302
rect 280 278 286 302
rect 222 222 226 278
rect 282 222 286 278
rect 222 209 228 222
rect 280 209 286 222
rect 222 198 286 209
rect 222 142 226 198
rect 282 142 286 198
rect 222 114 286 142
rect 316 519 380 825
rect 414 1196 478 1226
rect 414 1140 418 1196
rect 474 1140 478 1196
rect 414 1131 478 1140
rect 414 1116 420 1131
rect 472 1116 478 1131
rect 414 1060 418 1116
rect 474 1060 478 1116
rect 414 1036 420 1060
rect 472 1036 478 1060
rect 414 980 418 1036
rect 474 980 478 1036
rect 414 956 420 980
rect 472 956 478 980
rect 414 900 418 956
rect 474 900 478 956
rect 414 887 420 900
rect 472 887 478 900
rect 414 876 478 887
rect 414 820 418 876
rect 474 820 478 876
rect 414 792 478 820
rect 508 1197 572 1462
rect 508 1145 514 1197
rect 566 1145 572 1197
rect 508 1133 572 1145
rect 508 1081 514 1133
rect 566 1081 572 1133
rect 508 1069 572 1081
rect 508 1017 514 1069
rect 566 1017 572 1069
rect 508 1005 572 1017
rect 508 953 514 1005
rect 566 953 572 1005
rect 508 941 572 953
rect 508 889 514 941
rect 566 889 572 941
rect 508 877 572 889
rect 508 825 514 877
rect 566 825 572 877
rect 316 467 322 519
rect 374 467 380 519
rect 316 455 380 467
rect 316 403 322 455
rect 374 403 380 455
rect 316 391 380 403
rect 316 339 322 391
rect 374 339 380 391
rect 316 327 380 339
rect 316 275 322 327
rect 374 275 380 327
rect 316 263 380 275
rect 316 211 322 263
rect 374 211 380 263
rect 316 199 380 211
rect 316 147 322 199
rect 374 147 380 199
rect 316 114 380 147
rect 414 518 478 548
rect 414 462 418 518
rect 474 462 478 518
rect 414 453 478 462
rect 414 438 420 453
rect 472 438 478 453
rect 414 382 418 438
rect 474 382 478 438
rect 414 358 420 382
rect 472 358 478 382
rect 414 302 418 358
rect 474 302 478 358
rect 414 278 420 302
rect 472 278 478 302
rect 414 222 418 278
rect 474 222 478 278
rect 414 209 420 222
rect 472 209 478 222
rect 414 198 478 209
rect 414 142 418 198
rect 474 142 478 198
rect 414 114 478 142
rect 508 519 572 825
rect 606 1196 670 1226
rect 606 1140 610 1196
rect 666 1140 670 1196
rect 606 1131 670 1140
rect 606 1116 612 1131
rect 664 1116 670 1131
rect 606 1060 610 1116
rect 666 1060 670 1116
rect 606 1036 612 1060
rect 664 1036 670 1060
rect 606 980 610 1036
rect 666 980 670 1036
rect 606 956 612 980
rect 664 956 670 980
rect 606 900 610 956
rect 666 900 670 956
rect 606 887 612 900
rect 664 887 670 900
rect 606 876 670 887
rect 606 820 610 876
rect 666 820 670 876
rect 606 792 670 820
rect 700 1197 764 1462
rect 700 1145 706 1197
rect 758 1145 764 1197
rect 700 1133 764 1145
rect 700 1081 706 1133
rect 758 1081 764 1133
rect 700 1069 764 1081
rect 700 1017 706 1069
rect 758 1017 764 1069
rect 700 1005 764 1017
rect 700 953 706 1005
rect 758 953 764 1005
rect 700 941 764 953
rect 700 889 706 941
rect 758 889 764 941
rect 700 877 764 889
rect 700 825 706 877
rect 758 825 764 877
rect 508 467 514 519
rect 566 467 572 519
rect 508 455 572 467
rect 508 403 514 455
rect 566 403 572 455
rect 508 391 572 403
rect 508 339 514 391
rect 566 339 572 391
rect 508 327 572 339
rect 508 275 514 327
rect 566 275 572 327
rect 508 263 572 275
rect 508 211 514 263
rect 566 211 572 263
rect 508 199 572 211
rect 508 147 514 199
rect 566 147 572 199
rect 508 114 572 147
rect 606 518 670 548
rect 606 462 610 518
rect 666 462 670 518
rect 606 453 670 462
rect 606 438 612 453
rect 664 438 670 453
rect 606 382 610 438
rect 666 382 670 438
rect 606 358 612 382
rect 664 358 670 382
rect 606 302 610 358
rect 666 302 670 358
rect 606 278 612 302
rect 664 278 670 302
rect 606 222 610 278
rect 666 222 670 278
rect 606 209 612 222
rect 664 209 670 222
rect 606 198 670 209
rect 606 142 610 198
rect 666 142 670 198
rect 606 114 670 142
rect 700 519 764 825
rect 798 1196 862 1226
rect 798 1140 802 1196
rect 858 1140 862 1196
rect 798 1131 862 1140
rect 798 1116 804 1131
rect 856 1116 862 1131
rect 798 1060 802 1116
rect 858 1060 862 1116
rect 798 1036 804 1060
rect 856 1036 862 1060
rect 798 980 802 1036
rect 858 980 862 1036
rect 798 956 804 980
rect 856 956 862 980
rect 798 900 802 956
rect 858 900 862 956
rect 798 887 804 900
rect 856 887 862 900
rect 798 876 862 887
rect 798 820 802 876
rect 858 820 862 876
rect 798 792 862 820
rect 892 1197 956 1462
rect 892 1145 898 1197
rect 950 1145 956 1197
rect 892 1133 956 1145
rect 892 1081 898 1133
rect 950 1081 956 1133
rect 892 1069 956 1081
rect 892 1017 898 1069
rect 950 1017 956 1069
rect 892 1005 956 1017
rect 892 953 898 1005
rect 950 953 956 1005
rect 892 941 956 953
rect 892 889 898 941
rect 950 889 956 941
rect 892 877 956 889
rect 892 825 898 877
rect 950 825 956 877
rect 700 467 706 519
rect 758 467 764 519
rect 700 455 764 467
rect 700 403 706 455
rect 758 403 764 455
rect 700 391 764 403
rect 700 339 706 391
rect 758 339 764 391
rect 700 327 764 339
rect 700 275 706 327
rect 758 275 764 327
rect 700 263 764 275
rect 700 211 706 263
rect 758 211 764 263
rect 700 199 764 211
rect 700 147 706 199
rect 758 147 764 199
rect 700 114 764 147
rect 798 518 862 548
rect 798 462 802 518
rect 858 462 862 518
rect 798 453 862 462
rect 798 438 804 453
rect 856 438 862 453
rect 798 382 802 438
rect 858 382 862 438
rect 798 358 804 382
rect 856 358 862 382
rect 798 302 802 358
rect 858 302 862 358
rect 798 278 804 302
rect 856 278 862 302
rect 798 222 802 278
rect 858 222 862 278
rect 798 209 804 222
rect 856 209 862 222
rect 798 198 862 209
rect 798 142 802 198
rect 858 142 862 198
rect 798 114 862 142
rect 892 519 956 825
rect 990 1196 1054 1226
rect 990 1140 994 1196
rect 1050 1140 1054 1196
rect 990 1131 1054 1140
rect 990 1116 996 1131
rect 1048 1116 1054 1131
rect 990 1060 994 1116
rect 1050 1060 1054 1116
rect 990 1036 996 1060
rect 1048 1036 1054 1060
rect 990 980 994 1036
rect 1050 980 1054 1036
rect 990 956 996 980
rect 1048 956 1054 980
rect 990 900 994 956
rect 1050 900 1054 956
rect 990 887 996 900
rect 1048 887 1054 900
rect 990 876 1054 887
rect 990 820 994 876
rect 1050 820 1054 876
rect 990 792 1054 820
rect 1084 1197 1148 1462
rect 1084 1145 1090 1197
rect 1142 1145 1148 1197
rect 1084 1133 1148 1145
rect 1084 1081 1090 1133
rect 1142 1081 1148 1133
rect 1084 1069 1148 1081
rect 1084 1017 1090 1069
rect 1142 1017 1148 1069
rect 1084 1005 1148 1017
rect 1084 953 1090 1005
rect 1142 953 1148 1005
rect 1084 941 1148 953
rect 1084 889 1090 941
rect 1142 889 1148 941
rect 1084 877 1148 889
rect 1084 825 1090 877
rect 1142 825 1148 877
rect 892 467 898 519
rect 950 467 956 519
rect 892 455 956 467
rect 892 403 898 455
rect 950 403 956 455
rect 892 391 956 403
rect 892 339 898 391
rect 950 339 956 391
rect 892 327 956 339
rect 892 275 898 327
rect 950 275 956 327
rect 892 263 956 275
rect 892 211 898 263
rect 950 211 956 263
rect 892 199 956 211
rect 892 147 898 199
rect 950 147 956 199
rect 892 114 956 147
rect 990 518 1054 548
rect 990 462 994 518
rect 1050 462 1054 518
rect 990 453 1054 462
rect 990 438 996 453
rect 1048 438 1054 453
rect 990 382 994 438
rect 1050 382 1054 438
rect 990 358 996 382
rect 1048 358 1054 382
rect 990 302 994 358
rect 1050 302 1054 358
rect 990 278 996 302
rect 1048 278 1054 302
rect 990 222 994 278
rect 1050 222 1054 278
rect 990 209 996 222
rect 1048 209 1054 222
rect 990 198 1054 209
rect 990 142 994 198
rect 1050 142 1054 198
rect 990 114 1054 142
rect 1084 519 1148 825
rect 1182 1196 1246 1226
rect 1182 1140 1186 1196
rect 1242 1140 1246 1196
rect 1182 1131 1246 1140
rect 1182 1116 1188 1131
rect 1240 1116 1246 1131
rect 1182 1060 1186 1116
rect 1242 1060 1246 1116
rect 1182 1036 1188 1060
rect 1240 1036 1246 1060
rect 1182 980 1186 1036
rect 1242 980 1246 1036
rect 1182 956 1188 980
rect 1240 956 1246 980
rect 1182 900 1186 956
rect 1242 900 1246 956
rect 1182 887 1188 900
rect 1240 887 1246 900
rect 1182 876 1246 887
rect 1182 820 1186 876
rect 1242 820 1246 876
rect 1182 792 1246 820
rect 1276 1197 1340 1470
rect 1276 1145 1282 1197
rect 1334 1145 1340 1197
rect 1276 1133 1340 1145
rect 1276 1081 1282 1133
rect 1334 1081 1340 1133
rect 1276 1069 1340 1081
rect 1276 1017 1282 1069
rect 1334 1017 1340 1069
rect 1276 1005 1340 1017
rect 1276 953 1282 1005
rect 1334 953 1340 1005
rect 1276 941 1340 953
rect 1276 889 1282 941
rect 1334 889 1340 941
rect 1276 877 1340 889
rect 1276 825 1282 877
rect 1334 825 1340 877
rect 1084 467 1090 519
rect 1142 467 1148 519
rect 1084 455 1148 467
rect 1084 403 1090 455
rect 1142 403 1148 455
rect 1084 391 1148 403
rect 1084 339 1090 391
rect 1142 339 1148 391
rect 1084 327 1148 339
rect 1084 275 1090 327
rect 1142 275 1148 327
rect 1084 263 1148 275
rect 1084 211 1090 263
rect 1142 211 1148 263
rect 1084 199 1148 211
rect 1084 147 1090 199
rect 1142 147 1148 199
rect 1084 114 1148 147
rect 1182 518 1246 548
rect 1182 462 1186 518
rect 1242 462 1246 518
rect 1182 453 1246 462
rect 1182 438 1188 453
rect 1240 438 1246 453
rect 1182 382 1186 438
rect 1242 382 1246 438
rect 1182 358 1188 382
rect 1240 358 1246 382
rect 1182 302 1186 358
rect 1242 302 1246 358
rect 1182 278 1188 302
rect 1240 278 1246 302
rect 1182 222 1186 278
rect 1242 222 1246 278
rect 1182 209 1188 222
rect 1240 209 1246 222
rect 1182 198 1246 209
rect 1182 142 1186 198
rect 1242 142 1246 198
rect 1182 114 1246 142
rect 1276 519 1340 825
rect 1374 1196 1438 1226
rect 1374 1140 1378 1196
rect 1434 1140 1438 1196
rect 1374 1131 1438 1140
rect 1374 1116 1380 1131
rect 1432 1116 1438 1131
rect 1374 1060 1378 1116
rect 1434 1060 1438 1116
rect 1374 1036 1380 1060
rect 1432 1036 1438 1060
rect 1374 980 1378 1036
rect 1434 980 1438 1036
rect 1374 956 1380 980
rect 1432 956 1438 980
rect 1374 900 1378 956
rect 1434 900 1438 956
rect 1374 887 1380 900
rect 1432 887 1438 900
rect 1374 876 1438 887
rect 1374 820 1378 876
rect 1434 820 1438 876
rect 1374 792 1438 820
rect 1468 1197 1532 1470
rect 1468 1145 1474 1197
rect 1526 1145 1532 1197
rect 1468 1133 1532 1145
rect 1468 1081 1474 1133
rect 1526 1081 1532 1133
rect 1468 1069 1532 1081
rect 1468 1017 1474 1069
rect 1526 1017 1532 1069
rect 1468 1005 1532 1017
rect 1468 953 1474 1005
rect 1526 953 1532 1005
rect 1468 941 1532 953
rect 1468 889 1474 941
rect 1526 889 1532 941
rect 1468 877 1532 889
rect 1468 825 1474 877
rect 1526 825 1532 877
rect 1276 467 1282 519
rect 1334 467 1340 519
rect 1276 455 1340 467
rect 1276 403 1282 455
rect 1334 403 1340 455
rect 1276 391 1340 403
rect 1276 339 1282 391
rect 1334 339 1340 391
rect 1276 327 1340 339
rect 1276 275 1282 327
rect 1334 275 1340 327
rect 1276 263 1340 275
rect 1276 211 1282 263
rect 1334 211 1340 263
rect 1276 199 1340 211
rect 1276 147 1282 199
rect 1334 147 1340 199
rect 1276 114 1340 147
rect 1374 518 1438 548
rect 1374 462 1378 518
rect 1434 462 1438 518
rect 1374 453 1438 462
rect 1374 438 1380 453
rect 1432 438 1438 453
rect 1374 382 1378 438
rect 1434 382 1438 438
rect 1374 358 1380 382
rect 1432 358 1438 382
rect 1374 302 1378 358
rect 1434 302 1438 358
rect 1374 278 1380 302
rect 1432 278 1438 302
rect 1374 222 1378 278
rect 1434 222 1438 278
rect 1374 209 1380 222
rect 1432 209 1438 222
rect 1374 198 1438 209
rect 1374 142 1378 198
rect 1434 142 1438 198
rect 1374 114 1438 142
rect 1468 519 1532 825
rect 1566 1196 1630 1226
rect 1566 1140 1570 1196
rect 1626 1140 1630 1196
rect 1566 1131 1630 1140
rect 1566 1116 1572 1131
rect 1624 1116 1630 1131
rect 1566 1060 1570 1116
rect 1626 1060 1630 1116
rect 1566 1036 1572 1060
rect 1624 1036 1630 1060
rect 1566 980 1570 1036
rect 1626 980 1630 1036
rect 1566 956 1572 980
rect 1624 956 1630 980
rect 1566 900 1570 956
rect 1626 900 1630 956
rect 1566 887 1572 900
rect 1624 887 1630 900
rect 1566 876 1630 887
rect 1566 820 1570 876
rect 1626 820 1630 876
rect 1566 792 1630 820
rect 1660 1197 1724 1470
rect 1660 1145 1666 1197
rect 1718 1145 1724 1197
rect 1660 1133 1724 1145
rect 1660 1081 1666 1133
rect 1718 1081 1724 1133
rect 1660 1069 1724 1081
rect 1660 1017 1666 1069
rect 1718 1017 1724 1069
rect 1660 1005 1724 1017
rect 1660 953 1666 1005
rect 1718 953 1724 1005
rect 1660 941 1724 953
rect 1660 889 1666 941
rect 1718 889 1724 941
rect 1660 877 1724 889
rect 1660 825 1666 877
rect 1718 825 1724 877
rect 1468 467 1474 519
rect 1526 467 1532 519
rect 1468 455 1532 467
rect 1468 403 1474 455
rect 1526 403 1532 455
rect 1468 391 1532 403
rect 1468 339 1474 391
rect 1526 339 1532 391
rect 1468 327 1532 339
rect 1468 275 1474 327
rect 1526 275 1532 327
rect 1468 263 1532 275
rect 1468 211 1474 263
rect 1526 211 1532 263
rect 1468 199 1532 211
rect 1468 147 1474 199
rect 1526 147 1532 199
rect 1468 114 1532 147
rect 1566 518 1630 548
rect 1566 462 1570 518
rect 1626 462 1630 518
rect 1566 453 1630 462
rect 1566 438 1572 453
rect 1624 438 1630 453
rect 1566 382 1570 438
rect 1626 382 1630 438
rect 1566 358 1572 382
rect 1624 358 1630 382
rect 1566 302 1570 358
rect 1626 302 1630 358
rect 1566 278 1572 302
rect 1624 278 1630 302
rect 1566 222 1570 278
rect 1626 222 1630 278
rect 1566 209 1572 222
rect 1624 209 1630 222
rect 1566 198 1630 209
rect 1566 142 1570 198
rect 1626 142 1630 198
rect 1566 114 1630 142
rect 1660 519 1724 825
rect 1758 1196 1822 1226
rect 1758 1140 1762 1196
rect 1818 1140 1822 1196
rect 1758 1131 1822 1140
rect 1758 1116 1764 1131
rect 1816 1116 1822 1131
rect 1758 1060 1762 1116
rect 1818 1060 1822 1116
rect 1758 1036 1764 1060
rect 1816 1036 1822 1060
rect 1758 980 1762 1036
rect 1818 980 1822 1036
rect 1758 956 1764 980
rect 1816 956 1822 980
rect 1758 900 1762 956
rect 1818 900 1822 956
rect 1758 887 1764 900
rect 1816 887 1822 900
rect 1758 876 1822 887
rect 1758 820 1762 876
rect 1818 820 1822 876
rect 1758 792 1822 820
rect 1660 467 1666 519
rect 1718 467 1724 519
rect 1660 455 1724 467
rect 1660 403 1666 455
rect 1718 403 1724 455
rect 1660 391 1724 403
rect 1660 339 1666 391
rect 1718 339 1724 391
rect 1660 327 1724 339
rect 1660 275 1666 327
rect 1718 275 1724 327
rect 1660 263 1724 275
rect 1660 211 1666 263
rect 1718 211 1724 263
rect 1660 199 1724 211
rect 1660 147 1666 199
rect 1718 147 1724 199
rect 1660 114 1724 147
rect 1758 518 1822 548
rect 1758 462 1762 518
rect 1818 462 1822 518
rect 1758 453 1822 462
rect 1758 438 1764 453
rect 1816 438 1822 453
rect 1758 382 1762 438
rect 1818 382 1822 438
rect 1758 358 1764 382
rect 1816 358 1822 382
rect 1758 302 1762 358
rect 1818 302 1822 358
rect 1758 278 1764 302
rect 1816 278 1822 302
rect 1758 222 1762 278
rect 1818 222 1822 278
rect 1758 209 1764 222
rect 1816 209 1822 222
rect 1758 198 1822 209
rect 1758 142 1762 198
rect 1818 142 1822 198
rect 1758 114 1822 142
rect 34 -370 100 -342
rect 34 -426 38 -370
rect 94 -426 100 -370
rect 34 -432 40 -426
rect 92 -432 100 -426
rect 34 -444 100 -432
rect 34 -450 40 -444
rect 92 -450 100 -444
rect 34 -506 38 -450
rect 94 -506 100 -450
rect 34 -534 100 -506
rect 130 -379 194 -344
rect 130 -431 136 -379
rect 188 -431 194 -379
rect 130 -443 194 -431
rect 130 -495 136 -443
rect 188 -495 194 -443
rect 34 -778 100 -750
rect 34 -834 38 -778
rect 94 -834 100 -778
rect 34 -840 40 -834
rect 92 -840 100 -834
rect 34 -852 100 -840
rect 34 -858 40 -852
rect 92 -858 100 -852
rect 34 -914 38 -858
rect 94 -914 100 -858
rect 34 -942 100 -914
rect 130 -789 194 -495
rect 226 -370 292 -342
rect 226 -426 230 -370
rect 286 -426 292 -370
rect 226 -432 232 -426
rect 284 -432 292 -426
rect 226 -444 292 -432
rect 226 -450 232 -444
rect 284 -450 292 -444
rect 226 -506 230 -450
rect 286 -506 292 -450
rect 226 -534 292 -506
rect 322 -379 386 -344
rect 322 -431 328 -379
rect 380 -431 386 -379
rect 322 -443 386 -431
rect 322 -495 328 -443
rect 380 -495 386 -443
rect 130 -841 136 -789
rect 188 -841 194 -789
rect 130 -853 194 -841
rect 130 -905 136 -853
rect 188 -905 194 -853
rect 130 -1142 194 -905
rect 226 -778 292 -750
rect 226 -834 230 -778
rect 286 -834 292 -778
rect 226 -840 232 -834
rect 284 -840 292 -834
rect 226 -852 292 -840
rect 226 -858 232 -852
rect 284 -858 292 -852
rect 226 -914 230 -858
rect 286 -914 292 -858
rect 226 -942 292 -914
rect 322 -789 386 -495
rect 418 -370 484 -342
rect 418 -426 422 -370
rect 478 -426 484 -370
rect 418 -432 424 -426
rect 476 -432 484 -426
rect 418 -444 484 -432
rect 418 -450 424 -444
rect 476 -450 484 -444
rect 418 -506 422 -450
rect 478 -506 484 -450
rect 418 -534 484 -506
rect 514 -379 578 -344
rect 514 -431 520 -379
rect 572 -431 578 -379
rect 514 -443 578 -431
rect 514 -495 520 -443
rect 572 -495 578 -443
rect 322 -841 328 -789
rect 380 -841 386 -789
rect 322 -853 386 -841
rect 322 -905 328 -853
rect 380 -905 386 -853
rect 322 -1142 386 -905
rect 418 -778 484 -750
rect 418 -834 422 -778
rect 478 -834 484 -778
rect 418 -840 424 -834
rect 476 -840 484 -834
rect 418 -852 484 -840
rect 418 -858 424 -852
rect 476 -858 484 -852
rect 418 -914 422 -858
rect 478 -914 484 -858
rect 418 -942 484 -914
rect 514 -789 578 -495
rect 610 -370 676 -342
rect 610 -426 614 -370
rect 670 -426 676 -370
rect 610 -432 616 -426
rect 668 -432 676 -426
rect 610 -444 676 -432
rect 610 -450 616 -444
rect 668 -450 676 -444
rect 610 -506 614 -450
rect 670 -506 676 -450
rect 610 -534 676 -506
rect 706 -379 770 -344
rect 706 -431 712 -379
rect 764 -431 770 -379
rect 706 -443 770 -431
rect 706 -495 712 -443
rect 764 -495 770 -443
rect 514 -841 520 -789
rect 572 -841 578 -789
rect 514 -853 578 -841
rect 514 -905 520 -853
rect 572 -905 578 -853
rect 514 -1142 578 -905
rect 610 -778 676 -750
rect 610 -834 614 -778
rect 670 -834 676 -778
rect 610 -840 616 -834
rect 668 -840 676 -834
rect 610 -852 676 -840
rect 610 -858 616 -852
rect 668 -858 676 -852
rect 610 -914 614 -858
rect 670 -914 676 -858
rect 610 -942 676 -914
rect 706 -789 770 -495
rect 802 -370 868 -342
rect 802 -426 806 -370
rect 862 -426 868 -370
rect 802 -432 808 -426
rect 860 -432 868 -426
rect 802 -444 868 -432
rect 802 -450 808 -444
rect 860 -450 868 -444
rect 802 -506 806 -450
rect 862 -506 868 -450
rect 802 -534 868 -506
rect 898 -379 962 -344
rect 898 -431 904 -379
rect 956 -431 962 -379
rect 898 -443 962 -431
rect 898 -495 904 -443
rect 956 -495 962 -443
rect 706 -841 712 -789
rect 764 -841 770 -789
rect 706 -853 770 -841
rect 706 -905 712 -853
rect 764 -905 770 -853
rect 706 -1142 770 -905
rect 802 -778 868 -750
rect 802 -834 806 -778
rect 862 -834 868 -778
rect 802 -840 808 -834
rect 860 -840 868 -834
rect 802 -852 868 -840
rect 802 -858 808 -852
rect 860 -858 868 -852
rect 802 -914 806 -858
rect 862 -914 868 -858
rect 802 -942 868 -914
rect 898 -789 962 -495
rect 994 -370 1060 -342
rect 994 -426 998 -370
rect 1054 -426 1060 -370
rect 994 -432 1000 -426
rect 1052 -432 1060 -426
rect 994 -444 1060 -432
rect 994 -450 1000 -444
rect 1052 -450 1060 -444
rect 994 -506 998 -450
rect 1054 -506 1060 -450
rect 994 -534 1060 -506
rect 1090 -379 1154 -344
rect 1090 -431 1096 -379
rect 1148 -431 1154 -379
rect 1090 -443 1154 -431
rect 1090 -495 1096 -443
rect 1148 -495 1154 -443
rect 898 -841 904 -789
rect 956 -841 962 -789
rect 898 -853 962 -841
rect 898 -905 904 -853
rect 956 -905 962 -853
rect 898 -1142 962 -905
rect 994 -778 1060 -750
rect 994 -834 998 -778
rect 1054 -834 1060 -778
rect 994 -840 1000 -834
rect 1052 -840 1060 -834
rect 994 -852 1060 -840
rect 994 -858 1000 -852
rect 1052 -858 1060 -852
rect 994 -914 998 -858
rect 1054 -914 1060 -858
rect 994 -942 1060 -914
rect 1090 -789 1154 -495
rect 1186 -370 1252 -342
rect 1186 -426 1190 -370
rect 1246 -426 1252 -370
rect 1186 -432 1192 -426
rect 1244 -432 1252 -426
rect 1186 -444 1252 -432
rect 1186 -450 1192 -444
rect 1244 -450 1252 -444
rect 1186 -506 1190 -450
rect 1246 -506 1252 -450
rect 1186 -534 1252 -506
rect 1282 -379 1346 -344
rect 1282 -431 1288 -379
rect 1340 -431 1346 -379
rect 1282 -443 1346 -431
rect 1282 -495 1288 -443
rect 1340 -495 1346 -443
rect 1090 -841 1096 -789
rect 1148 -841 1154 -789
rect 1090 -853 1154 -841
rect 1090 -905 1096 -853
rect 1148 -905 1154 -853
rect 1090 -1142 1154 -905
rect 1186 -778 1252 -750
rect 1186 -834 1190 -778
rect 1246 -834 1252 -778
rect 1186 -840 1192 -834
rect 1244 -840 1252 -834
rect 1186 -852 1252 -840
rect 1186 -858 1192 -852
rect 1244 -858 1252 -852
rect 1186 -914 1190 -858
rect 1246 -914 1252 -858
rect 1186 -942 1252 -914
rect 1282 -789 1346 -495
rect 1378 -370 1444 -342
rect 1378 -426 1382 -370
rect 1438 -426 1444 -370
rect 1378 -432 1384 -426
rect 1436 -432 1444 -426
rect 1378 -444 1444 -432
rect 1378 -450 1384 -444
rect 1436 -450 1444 -444
rect 1378 -506 1382 -450
rect 1438 -506 1444 -450
rect 1378 -534 1444 -506
rect 1474 -379 1538 -344
rect 1474 -431 1480 -379
rect 1532 -431 1538 -379
rect 1474 -443 1538 -431
rect 1474 -495 1480 -443
rect 1532 -495 1538 -443
rect 1282 -841 1288 -789
rect 1340 -841 1346 -789
rect 1282 -853 1346 -841
rect 1282 -905 1288 -853
rect 1340 -905 1346 -853
rect 1282 -1142 1346 -905
rect 1378 -778 1444 -750
rect 1378 -834 1382 -778
rect 1438 -834 1444 -778
rect 1378 -840 1384 -834
rect 1436 -840 1444 -834
rect 1378 -852 1444 -840
rect 1378 -858 1384 -852
rect 1436 -858 1444 -852
rect 1378 -914 1382 -858
rect 1438 -914 1444 -858
rect 1378 -942 1444 -914
rect 1474 -789 1538 -495
rect 1570 -370 1636 -342
rect 1570 -426 1574 -370
rect 1630 -426 1636 -370
rect 1570 -432 1576 -426
rect 1628 -432 1636 -426
rect 1570 -444 1636 -432
rect 1570 -450 1576 -444
rect 1628 -450 1636 -444
rect 1570 -506 1574 -450
rect 1630 -506 1636 -450
rect 1570 -534 1636 -506
rect 1666 -379 1730 -344
rect 1666 -431 1672 -379
rect 1724 -431 1730 -379
rect 1666 -443 1730 -431
rect 1666 -495 1672 -443
rect 1724 -495 1730 -443
rect 1474 -841 1480 -789
rect 1532 -841 1538 -789
rect 1474 -853 1538 -841
rect 1474 -905 1480 -853
rect 1532 -905 1538 -853
rect 1474 -1142 1538 -905
rect 1570 -778 1636 -750
rect 1570 -834 1574 -778
rect 1630 -834 1636 -778
rect 1570 -840 1576 -834
rect 1628 -840 1636 -834
rect 1570 -852 1636 -840
rect 1570 -858 1576 -852
rect 1628 -858 1636 -852
rect 1570 -914 1574 -858
rect 1630 -914 1636 -858
rect 1570 -942 1636 -914
rect 1666 -789 1730 -495
rect 1762 -370 1828 -342
rect 1762 -426 1766 -370
rect 1822 -426 1828 -370
rect 1762 -432 1768 -426
rect 1820 -432 1828 -426
rect 1762 -444 1828 -432
rect 1762 -450 1768 -444
rect 1820 -450 1828 -444
rect 1762 -506 1766 -450
rect 1822 -506 1828 -450
rect 1762 -534 1828 -506
rect 1666 -841 1672 -789
rect 1724 -841 1730 -789
rect 1666 -853 1730 -841
rect 1666 -905 1672 -853
rect 1724 -905 1730 -853
rect 1666 -1142 1730 -905
rect 1762 -778 1828 -750
rect 1762 -834 1766 -778
rect 1822 -834 1828 -778
rect 1762 -840 1768 -834
rect 1820 -840 1828 -834
rect 1762 -852 1828 -840
rect 1762 -858 1768 -852
rect 1820 -858 1828 -852
rect 1762 -914 1766 -858
rect 1822 -914 1828 -858
rect 1762 -942 1828 -914
rect -84 -1164 1940 -1142
rect -104 -1168 1958 -1164
rect -104 -1220 -57 -1168
rect -5 -1220 7 -1168
rect 59 -1220 71 -1168
rect 123 -1220 135 -1168
rect 187 -1220 199 -1168
rect 251 -1220 263 -1168
rect 315 -1220 327 -1168
rect 379 -1220 391 -1168
rect 443 -1220 455 -1168
rect 507 -1220 519 -1168
rect 571 -1220 583 -1168
rect 635 -1220 647 -1168
rect 699 -1220 711 -1168
rect 763 -1220 775 -1168
rect 827 -1220 839 -1168
rect 891 -1220 903 -1168
rect 955 -1220 967 -1168
rect 1019 -1220 1031 -1168
rect 1083 -1220 1095 -1168
rect 1147 -1220 1159 -1168
rect 1211 -1220 1223 -1168
rect 1275 -1220 1287 -1168
rect 1339 -1220 1351 -1168
rect 1403 -1220 1415 -1168
rect 1467 -1220 1479 -1168
rect 1531 -1220 1543 -1168
rect 1595 -1220 1607 -1168
rect 1659 -1220 1671 -1168
rect 1723 -1220 1735 -1168
rect 1787 -1220 1799 -1168
rect 1851 -1220 1863 -1168
rect 1915 -1220 1958 -1168
rect -104 -1292 1958 -1220
<< via2 >>
rect 34 1195 90 1196
rect 34 1143 36 1195
rect 36 1143 88 1195
rect 88 1143 90 1195
rect 34 1140 90 1143
rect 34 1079 36 1116
rect 36 1079 88 1116
rect 88 1079 90 1116
rect 34 1067 90 1079
rect 34 1060 36 1067
rect 36 1060 88 1067
rect 88 1060 90 1067
rect 34 1015 36 1036
rect 36 1015 88 1036
rect 88 1015 90 1036
rect 34 1003 90 1015
rect 34 980 36 1003
rect 36 980 88 1003
rect 88 980 90 1003
rect 34 951 36 956
rect 36 951 88 956
rect 88 951 90 956
rect 34 939 90 951
rect 34 900 36 939
rect 36 900 88 939
rect 88 900 90 939
rect 34 875 90 876
rect 34 823 36 875
rect 36 823 88 875
rect 88 823 90 875
rect 34 820 90 823
rect 34 517 90 518
rect 34 465 36 517
rect 36 465 88 517
rect 88 465 90 517
rect 34 462 90 465
rect 34 401 36 438
rect 36 401 88 438
rect 88 401 90 438
rect 34 389 90 401
rect 34 382 36 389
rect 36 382 88 389
rect 88 382 90 389
rect 34 337 36 358
rect 36 337 88 358
rect 88 337 90 358
rect 34 325 90 337
rect 34 302 36 325
rect 36 302 88 325
rect 88 302 90 325
rect 34 273 36 278
rect 36 273 88 278
rect 88 273 90 278
rect 34 261 90 273
rect 34 222 36 261
rect 36 222 88 261
rect 88 222 90 261
rect 34 197 90 198
rect 34 145 36 197
rect 36 145 88 197
rect 88 145 90 197
rect 34 142 90 145
rect 226 1195 282 1196
rect 226 1143 228 1195
rect 228 1143 280 1195
rect 280 1143 282 1195
rect 226 1140 282 1143
rect 226 1079 228 1116
rect 228 1079 280 1116
rect 280 1079 282 1116
rect 226 1067 282 1079
rect 226 1060 228 1067
rect 228 1060 280 1067
rect 280 1060 282 1067
rect 226 1015 228 1036
rect 228 1015 280 1036
rect 280 1015 282 1036
rect 226 1003 282 1015
rect 226 980 228 1003
rect 228 980 280 1003
rect 280 980 282 1003
rect 226 951 228 956
rect 228 951 280 956
rect 280 951 282 956
rect 226 939 282 951
rect 226 900 228 939
rect 228 900 280 939
rect 280 900 282 939
rect 226 875 282 876
rect 226 823 228 875
rect 228 823 280 875
rect 280 823 282 875
rect 226 820 282 823
rect 226 517 282 518
rect 226 465 228 517
rect 228 465 280 517
rect 280 465 282 517
rect 226 462 282 465
rect 226 401 228 438
rect 228 401 280 438
rect 280 401 282 438
rect 226 389 282 401
rect 226 382 228 389
rect 228 382 280 389
rect 280 382 282 389
rect 226 337 228 358
rect 228 337 280 358
rect 280 337 282 358
rect 226 325 282 337
rect 226 302 228 325
rect 228 302 280 325
rect 280 302 282 325
rect 226 273 228 278
rect 228 273 280 278
rect 280 273 282 278
rect 226 261 282 273
rect 226 222 228 261
rect 228 222 280 261
rect 280 222 282 261
rect 226 197 282 198
rect 226 145 228 197
rect 228 145 280 197
rect 280 145 282 197
rect 226 142 282 145
rect 418 1195 474 1196
rect 418 1143 420 1195
rect 420 1143 472 1195
rect 472 1143 474 1195
rect 418 1140 474 1143
rect 418 1079 420 1116
rect 420 1079 472 1116
rect 472 1079 474 1116
rect 418 1067 474 1079
rect 418 1060 420 1067
rect 420 1060 472 1067
rect 472 1060 474 1067
rect 418 1015 420 1036
rect 420 1015 472 1036
rect 472 1015 474 1036
rect 418 1003 474 1015
rect 418 980 420 1003
rect 420 980 472 1003
rect 472 980 474 1003
rect 418 951 420 956
rect 420 951 472 956
rect 472 951 474 956
rect 418 939 474 951
rect 418 900 420 939
rect 420 900 472 939
rect 472 900 474 939
rect 418 875 474 876
rect 418 823 420 875
rect 420 823 472 875
rect 472 823 474 875
rect 418 820 474 823
rect 418 517 474 518
rect 418 465 420 517
rect 420 465 472 517
rect 472 465 474 517
rect 418 462 474 465
rect 418 401 420 438
rect 420 401 472 438
rect 472 401 474 438
rect 418 389 474 401
rect 418 382 420 389
rect 420 382 472 389
rect 472 382 474 389
rect 418 337 420 358
rect 420 337 472 358
rect 472 337 474 358
rect 418 325 474 337
rect 418 302 420 325
rect 420 302 472 325
rect 472 302 474 325
rect 418 273 420 278
rect 420 273 472 278
rect 472 273 474 278
rect 418 261 474 273
rect 418 222 420 261
rect 420 222 472 261
rect 472 222 474 261
rect 418 197 474 198
rect 418 145 420 197
rect 420 145 472 197
rect 472 145 474 197
rect 418 142 474 145
rect 610 1195 666 1196
rect 610 1143 612 1195
rect 612 1143 664 1195
rect 664 1143 666 1195
rect 610 1140 666 1143
rect 610 1079 612 1116
rect 612 1079 664 1116
rect 664 1079 666 1116
rect 610 1067 666 1079
rect 610 1060 612 1067
rect 612 1060 664 1067
rect 664 1060 666 1067
rect 610 1015 612 1036
rect 612 1015 664 1036
rect 664 1015 666 1036
rect 610 1003 666 1015
rect 610 980 612 1003
rect 612 980 664 1003
rect 664 980 666 1003
rect 610 951 612 956
rect 612 951 664 956
rect 664 951 666 956
rect 610 939 666 951
rect 610 900 612 939
rect 612 900 664 939
rect 664 900 666 939
rect 610 875 666 876
rect 610 823 612 875
rect 612 823 664 875
rect 664 823 666 875
rect 610 820 666 823
rect 610 517 666 518
rect 610 465 612 517
rect 612 465 664 517
rect 664 465 666 517
rect 610 462 666 465
rect 610 401 612 438
rect 612 401 664 438
rect 664 401 666 438
rect 610 389 666 401
rect 610 382 612 389
rect 612 382 664 389
rect 664 382 666 389
rect 610 337 612 358
rect 612 337 664 358
rect 664 337 666 358
rect 610 325 666 337
rect 610 302 612 325
rect 612 302 664 325
rect 664 302 666 325
rect 610 273 612 278
rect 612 273 664 278
rect 664 273 666 278
rect 610 261 666 273
rect 610 222 612 261
rect 612 222 664 261
rect 664 222 666 261
rect 610 197 666 198
rect 610 145 612 197
rect 612 145 664 197
rect 664 145 666 197
rect 610 142 666 145
rect 802 1195 858 1196
rect 802 1143 804 1195
rect 804 1143 856 1195
rect 856 1143 858 1195
rect 802 1140 858 1143
rect 802 1079 804 1116
rect 804 1079 856 1116
rect 856 1079 858 1116
rect 802 1067 858 1079
rect 802 1060 804 1067
rect 804 1060 856 1067
rect 856 1060 858 1067
rect 802 1015 804 1036
rect 804 1015 856 1036
rect 856 1015 858 1036
rect 802 1003 858 1015
rect 802 980 804 1003
rect 804 980 856 1003
rect 856 980 858 1003
rect 802 951 804 956
rect 804 951 856 956
rect 856 951 858 956
rect 802 939 858 951
rect 802 900 804 939
rect 804 900 856 939
rect 856 900 858 939
rect 802 875 858 876
rect 802 823 804 875
rect 804 823 856 875
rect 856 823 858 875
rect 802 820 858 823
rect 802 517 858 518
rect 802 465 804 517
rect 804 465 856 517
rect 856 465 858 517
rect 802 462 858 465
rect 802 401 804 438
rect 804 401 856 438
rect 856 401 858 438
rect 802 389 858 401
rect 802 382 804 389
rect 804 382 856 389
rect 856 382 858 389
rect 802 337 804 358
rect 804 337 856 358
rect 856 337 858 358
rect 802 325 858 337
rect 802 302 804 325
rect 804 302 856 325
rect 856 302 858 325
rect 802 273 804 278
rect 804 273 856 278
rect 856 273 858 278
rect 802 261 858 273
rect 802 222 804 261
rect 804 222 856 261
rect 856 222 858 261
rect 802 197 858 198
rect 802 145 804 197
rect 804 145 856 197
rect 856 145 858 197
rect 802 142 858 145
rect 994 1195 1050 1196
rect 994 1143 996 1195
rect 996 1143 1048 1195
rect 1048 1143 1050 1195
rect 994 1140 1050 1143
rect 994 1079 996 1116
rect 996 1079 1048 1116
rect 1048 1079 1050 1116
rect 994 1067 1050 1079
rect 994 1060 996 1067
rect 996 1060 1048 1067
rect 1048 1060 1050 1067
rect 994 1015 996 1036
rect 996 1015 1048 1036
rect 1048 1015 1050 1036
rect 994 1003 1050 1015
rect 994 980 996 1003
rect 996 980 1048 1003
rect 1048 980 1050 1003
rect 994 951 996 956
rect 996 951 1048 956
rect 1048 951 1050 956
rect 994 939 1050 951
rect 994 900 996 939
rect 996 900 1048 939
rect 1048 900 1050 939
rect 994 875 1050 876
rect 994 823 996 875
rect 996 823 1048 875
rect 1048 823 1050 875
rect 994 820 1050 823
rect 994 517 1050 518
rect 994 465 996 517
rect 996 465 1048 517
rect 1048 465 1050 517
rect 994 462 1050 465
rect 994 401 996 438
rect 996 401 1048 438
rect 1048 401 1050 438
rect 994 389 1050 401
rect 994 382 996 389
rect 996 382 1048 389
rect 1048 382 1050 389
rect 994 337 996 358
rect 996 337 1048 358
rect 1048 337 1050 358
rect 994 325 1050 337
rect 994 302 996 325
rect 996 302 1048 325
rect 1048 302 1050 325
rect 994 273 996 278
rect 996 273 1048 278
rect 1048 273 1050 278
rect 994 261 1050 273
rect 994 222 996 261
rect 996 222 1048 261
rect 1048 222 1050 261
rect 994 197 1050 198
rect 994 145 996 197
rect 996 145 1048 197
rect 1048 145 1050 197
rect 994 142 1050 145
rect 1186 1195 1242 1196
rect 1186 1143 1188 1195
rect 1188 1143 1240 1195
rect 1240 1143 1242 1195
rect 1186 1140 1242 1143
rect 1186 1079 1188 1116
rect 1188 1079 1240 1116
rect 1240 1079 1242 1116
rect 1186 1067 1242 1079
rect 1186 1060 1188 1067
rect 1188 1060 1240 1067
rect 1240 1060 1242 1067
rect 1186 1015 1188 1036
rect 1188 1015 1240 1036
rect 1240 1015 1242 1036
rect 1186 1003 1242 1015
rect 1186 980 1188 1003
rect 1188 980 1240 1003
rect 1240 980 1242 1003
rect 1186 951 1188 956
rect 1188 951 1240 956
rect 1240 951 1242 956
rect 1186 939 1242 951
rect 1186 900 1188 939
rect 1188 900 1240 939
rect 1240 900 1242 939
rect 1186 875 1242 876
rect 1186 823 1188 875
rect 1188 823 1240 875
rect 1240 823 1242 875
rect 1186 820 1242 823
rect 1186 517 1242 518
rect 1186 465 1188 517
rect 1188 465 1240 517
rect 1240 465 1242 517
rect 1186 462 1242 465
rect 1186 401 1188 438
rect 1188 401 1240 438
rect 1240 401 1242 438
rect 1186 389 1242 401
rect 1186 382 1188 389
rect 1188 382 1240 389
rect 1240 382 1242 389
rect 1186 337 1188 358
rect 1188 337 1240 358
rect 1240 337 1242 358
rect 1186 325 1242 337
rect 1186 302 1188 325
rect 1188 302 1240 325
rect 1240 302 1242 325
rect 1186 273 1188 278
rect 1188 273 1240 278
rect 1240 273 1242 278
rect 1186 261 1242 273
rect 1186 222 1188 261
rect 1188 222 1240 261
rect 1240 222 1242 261
rect 1186 197 1242 198
rect 1186 145 1188 197
rect 1188 145 1240 197
rect 1240 145 1242 197
rect 1186 142 1242 145
rect 1378 1195 1434 1196
rect 1378 1143 1380 1195
rect 1380 1143 1432 1195
rect 1432 1143 1434 1195
rect 1378 1140 1434 1143
rect 1378 1079 1380 1116
rect 1380 1079 1432 1116
rect 1432 1079 1434 1116
rect 1378 1067 1434 1079
rect 1378 1060 1380 1067
rect 1380 1060 1432 1067
rect 1432 1060 1434 1067
rect 1378 1015 1380 1036
rect 1380 1015 1432 1036
rect 1432 1015 1434 1036
rect 1378 1003 1434 1015
rect 1378 980 1380 1003
rect 1380 980 1432 1003
rect 1432 980 1434 1003
rect 1378 951 1380 956
rect 1380 951 1432 956
rect 1432 951 1434 956
rect 1378 939 1434 951
rect 1378 900 1380 939
rect 1380 900 1432 939
rect 1432 900 1434 939
rect 1378 875 1434 876
rect 1378 823 1380 875
rect 1380 823 1432 875
rect 1432 823 1434 875
rect 1378 820 1434 823
rect 1378 517 1434 518
rect 1378 465 1380 517
rect 1380 465 1432 517
rect 1432 465 1434 517
rect 1378 462 1434 465
rect 1378 401 1380 438
rect 1380 401 1432 438
rect 1432 401 1434 438
rect 1378 389 1434 401
rect 1378 382 1380 389
rect 1380 382 1432 389
rect 1432 382 1434 389
rect 1378 337 1380 358
rect 1380 337 1432 358
rect 1432 337 1434 358
rect 1378 325 1434 337
rect 1378 302 1380 325
rect 1380 302 1432 325
rect 1432 302 1434 325
rect 1378 273 1380 278
rect 1380 273 1432 278
rect 1432 273 1434 278
rect 1378 261 1434 273
rect 1378 222 1380 261
rect 1380 222 1432 261
rect 1432 222 1434 261
rect 1378 197 1434 198
rect 1378 145 1380 197
rect 1380 145 1432 197
rect 1432 145 1434 197
rect 1378 142 1434 145
rect 1570 1195 1626 1196
rect 1570 1143 1572 1195
rect 1572 1143 1624 1195
rect 1624 1143 1626 1195
rect 1570 1140 1626 1143
rect 1570 1079 1572 1116
rect 1572 1079 1624 1116
rect 1624 1079 1626 1116
rect 1570 1067 1626 1079
rect 1570 1060 1572 1067
rect 1572 1060 1624 1067
rect 1624 1060 1626 1067
rect 1570 1015 1572 1036
rect 1572 1015 1624 1036
rect 1624 1015 1626 1036
rect 1570 1003 1626 1015
rect 1570 980 1572 1003
rect 1572 980 1624 1003
rect 1624 980 1626 1003
rect 1570 951 1572 956
rect 1572 951 1624 956
rect 1624 951 1626 956
rect 1570 939 1626 951
rect 1570 900 1572 939
rect 1572 900 1624 939
rect 1624 900 1626 939
rect 1570 875 1626 876
rect 1570 823 1572 875
rect 1572 823 1624 875
rect 1624 823 1626 875
rect 1570 820 1626 823
rect 1570 517 1626 518
rect 1570 465 1572 517
rect 1572 465 1624 517
rect 1624 465 1626 517
rect 1570 462 1626 465
rect 1570 401 1572 438
rect 1572 401 1624 438
rect 1624 401 1626 438
rect 1570 389 1626 401
rect 1570 382 1572 389
rect 1572 382 1624 389
rect 1624 382 1626 389
rect 1570 337 1572 358
rect 1572 337 1624 358
rect 1624 337 1626 358
rect 1570 325 1626 337
rect 1570 302 1572 325
rect 1572 302 1624 325
rect 1624 302 1626 325
rect 1570 273 1572 278
rect 1572 273 1624 278
rect 1624 273 1626 278
rect 1570 261 1626 273
rect 1570 222 1572 261
rect 1572 222 1624 261
rect 1624 222 1626 261
rect 1570 197 1626 198
rect 1570 145 1572 197
rect 1572 145 1624 197
rect 1624 145 1626 197
rect 1570 142 1626 145
rect 1762 1195 1818 1196
rect 1762 1143 1764 1195
rect 1764 1143 1816 1195
rect 1816 1143 1818 1195
rect 1762 1140 1818 1143
rect 1762 1079 1764 1116
rect 1764 1079 1816 1116
rect 1816 1079 1818 1116
rect 1762 1067 1818 1079
rect 1762 1060 1764 1067
rect 1764 1060 1816 1067
rect 1816 1060 1818 1067
rect 1762 1015 1764 1036
rect 1764 1015 1816 1036
rect 1816 1015 1818 1036
rect 1762 1003 1818 1015
rect 1762 980 1764 1003
rect 1764 980 1816 1003
rect 1816 980 1818 1003
rect 1762 951 1764 956
rect 1764 951 1816 956
rect 1816 951 1818 956
rect 1762 939 1818 951
rect 1762 900 1764 939
rect 1764 900 1816 939
rect 1816 900 1818 939
rect 1762 875 1818 876
rect 1762 823 1764 875
rect 1764 823 1816 875
rect 1816 823 1818 875
rect 1762 820 1818 823
rect 1762 517 1818 518
rect 1762 465 1764 517
rect 1764 465 1816 517
rect 1816 465 1818 517
rect 1762 462 1818 465
rect 1762 401 1764 438
rect 1764 401 1816 438
rect 1816 401 1818 438
rect 1762 389 1818 401
rect 1762 382 1764 389
rect 1764 382 1816 389
rect 1816 382 1818 389
rect 1762 337 1764 358
rect 1764 337 1816 358
rect 1816 337 1818 358
rect 1762 325 1818 337
rect 1762 302 1764 325
rect 1764 302 1816 325
rect 1816 302 1818 325
rect 1762 273 1764 278
rect 1764 273 1816 278
rect 1816 273 1818 278
rect 1762 261 1818 273
rect 1762 222 1764 261
rect 1764 222 1816 261
rect 1816 222 1818 261
rect 1762 197 1818 198
rect 1762 145 1764 197
rect 1764 145 1816 197
rect 1816 145 1818 197
rect 1762 142 1818 145
rect 38 -380 94 -370
rect 38 -426 40 -380
rect 40 -426 92 -380
rect 92 -426 94 -380
rect 38 -496 40 -450
rect 40 -496 92 -450
rect 92 -496 94 -450
rect 38 -506 94 -496
rect 38 -788 94 -778
rect 38 -834 40 -788
rect 40 -834 92 -788
rect 92 -834 94 -788
rect 38 -904 40 -858
rect 40 -904 92 -858
rect 92 -904 94 -858
rect 38 -914 94 -904
rect 230 -380 286 -370
rect 230 -426 232 -380
rect 232 -426 284 -380
rect 284 -426 286 -380
rect 230 -496 232 -450
rect 232 -496 284 -450
rect 284 -496 286 -450
rect 230 -506 286 -496
rect 230 -788 286 -778
rect 230 -834 232 -788
rect 232 -834 284 -788
rect 284 -834 286 -788
rect 230 -904 232 -858
rect 232 -904 284 -858
rect 284 -904 286 -858
rect 230 -914 286 -904
rect 422 -380 478 -370
rect 422 -426 424 -380
rect 424 -426 476 -380
rect 476 -426 478 -380
rect 422 -496 424 -450
rect 424 -496 476 -450
rect 476 -496 478 -450
rect 422 -506 478 -496
rect 422 -788 478 -778
rect 422 -834 424 -788
rect 424 -834 476 -788
rect 476 -834 478 -788
rect 422 -904 424 -858
rect 424 -904 476 -858
rect 476 -904 478 -858
rect 422 -914 478 -904
rect 614 -380 670 -370
rect 614 -426 616 -380
rect 616 -426 668 -380
rect 668 -426 670 -380
rect 614 -496 616 -450
rect 616 -496 668 -450
rect 668 -496 670 -450
rect 614 -506 670 -496
rect 614 -788 670 -778
rect 614 -834 616 -788
rect 616 -834 668 -788
rect 668 -834 670 -788
rect 614 -904 616 -858
rect 616 -904 668 -858
rect 668 -904 670 -858
rect 614 -914 670 -904
rect 806 -380 862 -370
rect 806 -426 808 -380
rect 808 -426 860 -380
rect 860 -426 862 -380
rect 806 -496 808 -450
rect 808 -496 860 -450
rect 860 -496 862 -450
rect 806 -506 862 -496
rect 806 -788 862 -778
rect 806 -834 808 -788
rect 808 -834 860 -788
rect 860 -834 862 -788
rect 806 -904 808 -858
rect 808 -904 860 -858
rect 860 -904 862 -858
rect 806 -914 862 -904
rect 998 -380 1054 -370
rect 998 -426 1000 -380
rect 1000 -426 1052 -380
rect 1052 -426 1054 -380
rect 998 -496 1000 -450
rect 1000 -496 1052 -450
rect 1052 -496 1054 -450
rect 998 -506 1054 -496
rect 998 -788 1054 -778
rect 998 -834 1000 -788
rect 1000 -834 1052 -788
rect 1052 -834 1054 -788
rect 998 -904 1000 -858
rect 1000 -904 1052 -858
rect 1052 -904 1054 -858
rect 998 -914 1054 -904
rect 1190 -380 1246 -370
rect 1190 -426 1192 -380
rect 1192 -426 1244 -380
rect 1244 -426 1246 -380
rect 1190 -496 1192 -450
rect 1192 -496 1244 -450
rect 1244 -496 1246 -450
rect 1190 -506 1246 -496
rect 1190 -788 1246 -778
rect 1190 -834 1192 -788
rect 1192 -834 1244 -788
rect 1244 -834 1246 -788
rect 1190 -904 1192 -858
rect 1192 -904 1244 -858
rect 1244 -904 1246 -858
rect 1190 -914 1246 -904
rect 1382 -380 1438 -370
rect 1382 -426 1384 -380
rect 1384 -426 1436 -380
rect 1436 -426 1438 -380
rect 1382 -496 1384 -450
rect 1384 -496 1436 -450
rect 1436 -496 1438 -450
rect 1382 -506 1438 -496
rect 1382 -788 1438 -778
rect 1382 -834 1384 -788
rect 1384 -834 1436 -788
rect 1436 -834 1438 -788
rect 1382 -904 1384 -858
rect 1384 -904 1436 -858
rect 1436 -904 1438 -858
rect 1382 -914 1438 -904
rect 1574 -380 1630 -370
rect 1574 -426 1576 -380
rect 1576 -426 1628 -380
rect 1628 -426 1630 -380
rect 1574 -496 1576 -450
rect 1576 -496 1628 -450
rect 1628 -496 1630 -450
rect 1574 -506 1630 -496
rect 1574 -788 1630 -778
rect 1574 -834 1576 -788
rect 1576 -834 1628 -788
rect 1628 -834 1630 -788
rect 1574 -904 1576 -858
rect 1576 -904 1628 -858
rect 1628 -904 1630 -858
rect 1574 -914 1630 -904
rect 1766 -380 1822 -370
rect 1766 -426 1768 -380
rect 1768 -426 1820 -380
rect 1820 -426 1822 -380
rect 1766 -496 1768 -450
rect 1768 -496 1820 -450
rect 1820 -496 1822 -450
rect 1766 -506 1822 -496
rect 1766 -788 1822 -778
rect 1766 -834 1768 -788
rect 1768 -834 1820 -788
rect 1820 -834 1822 -788
rect 1766 -904 1768 -858
rect 1768 -904 1820 -858
rect 1820 -904 1822 -858
rect 1766 -914 1822 -904
<< metal3 >>
rect 28 1196 96 1228
rect 28 1140 34 1196
rect 90 1140 96 1196
rect 28 1116 96 1140
rect 28 1060 34 1116
rect 90 1060 96 1116
rect 28 1036 96 1060
rect 28 980 34 1036
rect 90 980 96 1036
rect 28 956 96 980
rect 28 900 34 956
rect 90 900 96 956
rect 28 876 96 900
rect 28 820 34 876
rect 90 820 96 876
rect 28 518 96 820
rect 28 462 34 518
rect 90 462 96 518
rect 28 438 96 462
rect 28 382 34 438
rect 90 382 96 438
rect 28 358 96 382
rect 28 302 34 358
rect 90 302 96 358
rect 28 278 96 302
rect 28 222 34 278
rect 90 222 96 278
rect 28 198 96 222
rect 28 142 34 198
rect 90 142 96 198
rect 28 -36 96 142
rect 220 1196 288 1228
rect 220 1140 226 1196
rect 282 1140 288 1196
rect 220 1116 288 1140
rect 220 1060 226 1116
rect 282 1060 288 1116
rect 220 1036 288 1060
rect 220 980 226 1036
rect 282 980 288 1036
rect 220 956 288 980
rect 220 900 226 956
rect 282 900 288 956
rect 220 876 288 900
rect 220 820 226 876
rect 282 820 288 876
rect 220 518 288 820
rect 220 462 226 518
rect 282 462 288 518
rect 220 438 288 462
rect 220 382 226 438
rect 282 382 288 438
rect 220 358 288 382
rect 220 302 226 358
rect 282 302 288 358
rect 220 278 288 302
rect 220 222 226 278
rect 282 222 288 278
rect 220 198 288 222
rect 220 142 226 198
rect 282 142 288 198
rect 220 -36 288 142
rect 412 1196 480 1228
rect 412 1140 418 1196
rect 474 1140 480 1196
rect 412 1116 480 1140
rect 412 1060 418 1116
rect 474 1060 480 1116
rect 412 1036 480 1060
rect 412 980 418 1036
rect 474 980 480 1036
rect 412 956 480 980
rect 412 900 418 956
rect 474 900 480 956
rect 412 876 480 900
rect 412 820 418 876
rect 474 820 480 876
rect 412 518 480 820
rect 412 462 418 518
rect 474 462 480 518
rect 412 438 480 462
rect 412 382 418 438
rect 474 382 480 438
rect 412 358 480 382
rect 412 302 418 358
rect 474 302 480 358
rect 412 278 480 302
rect 412 222 418 278
rect 474 222 480 278
rect 412 198 480 222
rect 412 142 418 198
rect 474 142 480 198
rect 412 -36 480 142
rect 604 1196 672 1228
rect 604 1140 610 1196
rect 666 1140 672 1196
rect 604 1116 672 1140
rect 604 1060 610 1116
rect 666 1060 672 1116
rect 604 1036 672 1060
rect 604 980 610 1036
rect 666 980 672 1036
rect 604 956 672 980
rect 604 900 610 956
rect 666 900 672 956
rect 604 876 672 900
rect 604 820 610 876
rect 666 820 672 876
rect 604 518 672 820
rect 604 462 610 518
rect 666 462 672 518
rect 604 438 672 462
rect 604 382 610 438
rect 666 382 672 438
rect 604 358 672 382
rect 604 302 610 358
rect 666 302 672 358
rect 604 278 672 302
rect 604 222 610 278
rect 666 222 672 278
rect 604 198 672 222
rect 604 142 610 198
rect 666 142 672 198
rect 604 -36 672 142
rect 796 1196 864 1228
rect 796 1140 802 1196
rect 858 1140 864 1196
rect 796 1116 864 1140
rect 796 1060 802 1116
rect 858 1060 864 1116
rect 796 1036 864 1060
rect 796 980 802 1036
rect 858 980 864 1036
rect 796 956 864 980
rect 796 900 802 956
rect 858 900 864 956
rect 796 876 864 900
rect 796 820 802 876
rect 858 820 864 876
rect 796 518 864 820
rect 796 462 802 518
rect 858 462 864 518
rect 796 438 864 462
rect 796 382 802 438
rect 858 382 864 438
rect 796 358 864 382
rect 796 302 802 358
rect 858 302 864 358
rect 796 278 864 302
rect 796 222 802 278
rect 858 222 864 278
rect 796 198 864 222
rect 796 142 802 198
rect 858 142 864 198
rect 796 -36 864 142
rect 988 1196 1056 1228
rect 988 1140 994 1196
rect 1050 1140 1056 1196
rect 988 1116 1056 1140
rect 988 1060 994 1116
rect 1050 1060 1056 1116
rect 988 1036 1056 1060
rect 988 980 994 1036
rect 1050 980 1056 1036
rect 988 956 1056 980
rect 988 900 994 956
rect 1050 900 1056 956
rect 988 876 1056 900
rect 988 820 994 876
rect 1050 820 1056 876
rect 988 518 1056 820
rect 988 462 994 518
rect 1050 462 1056 518
rect 988 438 1056 462
rect 988 382 994 438
rect 1050 382 1056 438
rect 988 358 1056 382
rect 988 302 994 358
rect 1050 302 1056 358
rect 988 278 1056 302
rect 988 222 994 278
rect 1050 222 1056 278
rect 988 198 1056 222
rect 988 142 994 198
rect 1050 142 1056 198
rect 988 -36 1056 142
rect 1180 1196 1248 1228
rect 1180 1140 1186 1196
rect 1242 1140 1248 1196
rect 1180 1116 1248 1140
rect 1180 1060 1186 1116
rect 1242 1060 1248 1116
rect 1180 1036 1248 1060
rect 1180 980 1186 1036
rect 1242 980 1248 1036
rect 1180 956 1248 980
rect 1180 900 1186 956
rect 1242 900 1248 956
rect 1180 876 1248 900
rect 1180 820 1186 876
rect 1242 820 1248 876
rect 1180 518 1248 820
rect 1180 462 1186 518
rect 1242 462 1248 518
rect 1180 438 1248 462
rect 1180 382 1186 438
rect 1242 382 1248 438
rect 1180 358 1248 382
rect 1180 302 1186 358
rect 1242 302 1248 358
rect 1180 278 1248 302
rect 1180 222 1186 278
rect 1242 222 1248 278
rect 1180 198 1248 222
rect 1180 142 1186 198
rect 1242 142 1248 198
rect 1180 -36 1248 142
rect 1372 1196 1440 1228
rect 1372 1140 1378 1196
rect 1434 1140 1440 1196
rect 1372 1116 1440 1140
rect 1372 1060 1378 1116
rect 1434 1060 1440 1116
rect 1372 1036 1440 1060
rect 1372 980 1378 1036
rect 1434 980 1440 1036
rect 1372 956 1440 980
rect 1372 900 1378 956
rect 1434 900 1440 956
rect 1372 876 1440 900
rect 1372 820 1378 876
rect 1434 820 1440 876
rect 1372 518 1440 820
rect 1372 462 1378 518
rect 1434 462 1440 518
rect 1372 438 1440 462
rect 1372 382 1378 438
rect 1434 382 1440 438
rect 1372 358 1440 382
rect 1372 302 1378 358
rect 1434 302 1440 358
rect 1372 278 1440 302
rect 1372 222 1378 278
rect 1434 222 1440 278
rect 1372 198 1440 222
rect 1372 142 1378 198
rect 1434 142 1440 198
rect 1372 -36 1440 142
rect 1564 1196 1632 1228
rect 1564 1140 1570 1196
rect 1626 1140 1632 1196
rect 1564 1116 1632 1140
rect 1564 1060 1570 1116
rect 1626 1060 1632 1116
rect 1564 1036 1632 1060
rect 1564 980 1570 1036
rect 1626 980 1632 1036
rect 1564 956 1632 980
rect 1564 900 1570 956
rect 1626 900 1632 956
rect 1564 876 1632 900
rect 1564 820 1570 876
rect 1626 820 1632 876
rect 1564 518 1632 820
rect 1564 462 1570 518
rect 1626 462 1632 518
rect 1564 438 1632 462
rect 1564 382 1570 438
rect 1626 382 1632 438
rect 1564 358 1632 382
rect 1564 302 1570 358
rect 1626 302 1632 358
rect 1564 278 1632 302
rect 1564 222 1570 278
rect 1626 222 1632 278
rect 1564 198 1632 222
rect 1564 142 1570 198
rect 1626 142 1632 198
rect 1564 -36 1632 142
rect 1756 1196 1824 1228
rect 1756 1140 1762 1196
rect 1818 1140 1824 1196
rect 1756 1116 1824 1140
rect 1756 1060 1762 1116
rect 1818 1060 1824 1116
rect 1756 1036 1824 1060
rect 1756 980 1762 1036
rect 1818 980 1824 1036
rect 1756 956 1824 980
rect 1756 900 1762 956
rect 1818 900 1824 956
rect 1756 876 1824 900
rect 1756 820 1762 876
rect 1818 820 1824 876
rect 1756 518 1824 820
rect 1756 462 1762 518
rect 1818 462 1824 518
rect 1756 438 1824 462
rect 1756 382 1762 438
rect 1818 382 1824 438
rect 1756 358 1824 382
rect 1756 302 1762 358
rect 1818 302 1824 358
rect 1756 278 1824 302
rect 1756 222 1762 278
rect 1818 222 1824 278
rect 1756 198 1824 222
rect 1756 142 1762 198
rect 1818 142 1824 198
rect 1756 -36 1824 142
rect 28 -200 1986 -36
rect 32 -370 100 -200
rect 32 -426 38 -370
rect 94 -426 100 -370
rect 32 -450 100 -426
rect 32 -506 38 -450
rect 94 -506 100 -450
rect 32 -778 100 -506
rect 32 -834 38 -778
rect 94 -834 100 -778
rect 32 -858 100 -834
rect 32 -914 38 -858
rect 94 -914 100 -858
rect 32 -942 100 -914
rect 224 -370 292 -200
rect 224 -426 230 -370
rect 286 -426 292 -370
rect 224 -450 292 -426
rect 224 -506 230 -450
rect 286 -506 292 -450
rect 224 -778 292 -506
rect 224 -834 230 -778
rect 286 -834 292 -778
rect 224 -858 292 -834
rect 224 -914 230 -858
rect 286 -914 292 -858
rect 224 -942 292 -914
rect 416 -370 484 -200
rect 416 -426 422 -370
rect 478 -426 484 -370
rect 416 -450 484 -426
rect 416 -506 422 -450
rect 478 -506 484 -450
rect 416 -778 484 -506
rect 416 -834 422 -778
rect 478 -834 484 -778
rect 416 -858 484 -834
rect 416 -914 422 -858
rect 478 -914 484 -858
rect 416 -942 484 -914
rect 608 -370 676 -200
rect 608 -426 614 -370
rect 670 -426 676 -370
rect 608 -450 676 -426
rect 608 -506 614 -450
rect 670 -506 676 -450
rect 608 -778 676 -506
rect 608 -834 614 -778
rect 670 -834 676 -778
rect 608 -858 676 -834
rect 608 -914 614 -858
rect 670 -914 676 -858
rect 608 -942 676 -914
rect 800 -370 868 -200
rect 800 -426 806 -370
rect 862 -426 868 -370
rect 800 -450 868 -426
rect 800 -506 806 -450
rect 862 -506 868 -450
rect 800 -778 868 -506
rect 800 -834 806 -778
rect 862 -834 868 -778
rect 800 -858 868 -834
rect 800 -914 806 -858
rect 862 -914 868 -858
rect 800 -942 868 -914
rect 992 -370 1060 -200
rect 992 -426 998 -370
rect 1054 -426 1060 -370
rect 992 -450 1060 -426
rect 992 -506 998 -450
rect 1054 -506 1060 -450
rect 992 -778 1060 -506
rect 992 -834 998 -778
rect 1054 -834 1060 -778
rect 992 -858 1060 -834
rect 992 -914 998 -858
rect 1054 -914 1060 -858
rect 992 -942 1060 -914
rect 1184 -370 1252 -200
rect 1184 -426 1190 -370
rect 1246 -426 1252 -370
rect 1184 -450 1252 -426
rect 1184 -506 1190 -450
rect 1246 -506 1252 -450
rect 1184 -778 1252 -506
rect 1184 -834 1190 -778
rect 1246 -834 1252 -778
rect 1184 -858 1252 -834
rect 1184 -914 1190 -858
rect 1246 -914 1252 -858
rect 1184 -942 1252 -914
rect 1376 -370 1444 -200
rect 1376 -426 1382 -370
rect 1438 -426 1444 -370
rect 1376 -450 1444 -426
rect 1376 -506 1382 -450
rect 1438 -506 1444 -450
rect 1376 -778 1444 -506
rect 1376 -834 1382 -778
rect 1438 -834 1444 -778
rect 1376 -858 1444 -834
rect 1376 -914 1382 -858
rect 1438 -914 1444 -858
rect 1376 -942 1444 -914
rect 1568 -370 1636 -200
rect 1568 -426 1574 -370
rect 1630 -426 1636 -370
rect 1568 -450 1636 -426
rect 1568 -506 1574 -450
rect 1630 -506 1636 -450
rect 1568 -778 1636 -506
rect 1568 -834 1574 -778
rect 1630 -834 1636 -778
rect 1568 -858 1636 -834
rect 1568 -914 1574 -858
rect 1630 -914 1636 -858
rect 1568 -942 1636 -914
rect 1760 -370 1828 -200
rect 1760 -426 1766 -370
rect 1822 -426 1828 -370
rect 1760 -450 1828 -426
rect 1760 -506 1766 -450
rect 1822 -506 1828 -450
rect 1760 -778 1828 -506
rect 1760 -834 1766 -778
rect 1822 -834 1828 -778
rect 1760 -858 1828 -834
rect 1760 -914 1766 -858
rect 1822 -914 1828 -858
rect 1760 -942 1828 -914
use sky130_fd_pr__nfet_01v8_BBTBMZ  sky130_fd_pr__nfet_01v8_BBTBMZ_0
timestamp 1627926120
transform 1 0 929 0 1 -641
box -995 -475 995 475
use sky130_fd_pr__pfet_01v8_VNEHM9  sky130_fd_pr__pfet_01v8_VNEHM9_0
timestamp 1627926120
transform 1 0 925 0 1 673
box -1031 -779 1031 779
<< labels >>
rlabel metal2 s -94 -1278 1952 -1176 4 GND
port 1 nsew
rlabel metal3 s 1934 -200 1986 -36 4 out
port 2 nsew
rlabel metal2 s -100 1480 1946 1582 4 VDD
port 3 nsew
rlabel metal1 s -160 -220 -16 -16 4 in
port 4 nsew
<< end >>
