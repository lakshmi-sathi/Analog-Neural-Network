magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_p >>
rect -1901 381 -1843 387
rect -1709 381 -1651 387
rect -1517 381 -1459 387
rect -1325 381 -1267 387
rect -1133 381 -1075 387
rect -941 381 -883 387
rect -749 381 -691 387
rect -557 381 -499 387
rect -365 381 -307 387
rect -173 381 -115 387
rect 19 381 77 387
rect 211 381 269 387
rect 403 381 461 387
rect 595 381 653 387
rect 787 381 845 387
rect 979 381 1037 387
rect 1171 381 1229 387
rect 1363 381 1421 387
rect 1555 381 1613 387
rect 1747 381 1805 387
rect 1939 381 1997 387
rect -1901 347 -1889 381
rect -1709 347 -1697 381
rect -1517 347 -1505 381
rect -1325 347 -1313 381
rect -1133 347 -1121 381
rect -941 347 -929 381
rect -749 347 -737 381
rect -557 347 -545 381
rect -365 347 -353 381
rect -173 347 -161 381
rect 19 347 31 381
rect 211 347 223 381
rect 403 347 415 381
rect 595 347 607 381
rect 787 347 799 381
rect 979 347 991 381
rect 1171 347 1183 381
rect 1363 347 1375 381
rect 1555 347 1567 381
rect 1747 347 1759 381
rect 1939 347 1951 381
rect -1901 341 -1843 347
rect -1709 341 -1651 347
rect -1517 341 -1459 347
rect -1325 341 -1267 347
rect -1133 341 -1075 347
rect -941 341 -883 347
rect -749 341 -691 347
rect -557 341 -499 347
rect -365 341 -307 347
rect -173 341 -115 347
rect 19 341 77 347
rect 211 341 269 347
rect 403 341 461 347
rect 595 341 653 347
rect 787 341 845 347
rect 979 341 1037 347
rect 1171 341 1229 347
rect 1363 341 1421 347
rect 1555 341 1613 347
rect 1747 341 1805 347
rect 1939 341 1997 347
rect -1997 -347 -1939 -341
rect -1805 -347 -1747 -341
rect -1613 -347 -1555 -341
rect -1421 -347 -1363 -341
rect -1229 -347 -1171 -341
rect -1037 -347 -979 -341
rect -845 -347 -787 -341
rect -653 -347 -595 -341
rect -461 -347 -403 -341
rect -269 -347 -211 -341
rect -77 -347 -19 -341
rect 115 -347 173 -341
rect 307 -347 365 -341
rect 499 -347 557 -341
rect 691 -347 749 -341
rect 883 -347 941 -341
rect 1075 -347 1133 -341
rect 1267 -347 1325 -341
rect 1459 -347 1517 -341
rect 1651 -347 1709 -341
rect 1843 -347 1901 -341
rect -1997 -381 -1985 -347
rect -1805 -381 -1793 -347
rect -1613 -381 -1601 -347
rect -1421 -381 -1409 -347
rect -1229 -381 -1217 -347
rect -1037 -381 -1025 -347
rect -845 -381 -833 -347
rect -653 -381 -641 -347
rect -461 -381 -449 -347
rect -269 -381 -257 -347
rect -77 -381 -65 -347
rect 115 -381 127 -347
rect 307 -381 319 -347
rect 499 -381 511 -347
rect 691 -381 703 -347
rect 883 -381 895 -347
rect 1075 -381 1087 -347
rect 1267 -381 1279 -347
rect 1459 -381 1471 -347
rect 1651 -381 1663 -347
rect 1843 -381 1855 -347
rect -1997 -387 -1939 -381
rect -1805 -387 -1747 -381
rect -1613 -387 -1555 -381
rect -1421 -387 -1363 -381
rect -1229 -387 -1171 -381
rect -1037 -387 -979 -381
rect -845 -387 -787 -381
rect -653 -387 -595 -381
rect -461 -387 -403 -381
rect -269 -387 -211 -381
rect -77 -387 -19 -381
rect 115 -387 173 -381
rect 307 -387 365 -381
rect 499 -387 557 -381
rect 691 -387 749 -381
rect 883 -387 941 -381
rect 1075 -387 1133 -381
rect 1267 -387 1325 -381
rect 1459 -387 1517 -381
rect 1651 -387 1709 -381
rect 1843 -387 1901 -381
<< nwell >>
rect -1985 362 2081 400
rect -2081 -362 2081 362
rect -2081 -400 1985 -362
<< pmos >>
rect -1983 -300 -1953 300
rect -1887 -300 -1857 300
rect -1791 -300 -1761 300
rect -1695 -300 -1665 300
rect -1599 -300 -1569 300
rect -1503 -300 -1473 300
rect -1407 -300 -1377 300
rect -1311 -300 -1281 300
rect -1215 -300 -1185 300
rect -1119 -300 -1089 300
rect -1023 -300 -993 300
rect -927 -300 -897 300
rect -831 -300 -801 300
rect -735 -300 -705 300
rect -639 -300 -609 300
rect -543 -300 -513 300
rect -447 -300 -417 300
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
rect 417 -300 447 300
rect 513 -300 543 300
rect 609 -300 639 300
rect 705 -300 735 300
rect 801 -300 831 300
rect 897 -300 927 300
rect 993 -300 1023 300
rect 1089 -300 1119 300
rect 1185 -300 1215 300
rect 1281 -300 1311 300
rect 1377 -300 1407 300
rect 1473 -300 1503 300
rect 1569 -300 1599 300
rect 1665 -300 1695 300
rect 1761 -300 1791 300
rect 1857 -300 1887 300
rect 1953 -300 1983 300
<< pdiff >>
rect -2045 255 -1983 300
rect -2045 221 -2033 255
rect -1999 221 -1983 255
rect -2045 187 -1983 221
rect -2045 153 -2033 187
rect -1999 153 -1983 187
rect -2045 119 -1983 153
rect -2045 85 -2033 119
rect -1999 85 -1983 119
rect -2045 51 -1983 85
rect -2045 17 -2033 51
rect -1999 17 -1983 51
rect -2045 -17 -1983 17
rect -2045 -51 -2033 -17
rect -1999 -51 -1983 -17
rect -2045 -85 -1983 -51
rect -2045 -119 -2033 -85
rect -1999 -119 -1983 -85
rect -2045 -153 -1983 -119
rect -2045 -187 -2033 -153
rect -1999 -187 -1983 -153
rect -2045 -221 -1983 -187
rect -2045 -255 -2033 -221
rect -1999 -255 -1983 -221
rect -2045 -300 -1983 -255
rect -1953 255 -1887 300
rect -1953 221 -1937 255
rect -1903 221 -1887 255
rect -1953 187 -1887 221
rect -1953 153 -1937 187
rect -1903 153 -1887 187
rect -1953 119 -1887 153
rect -1953 85 -1937 119
rect -1903 85 -1887 119
rect -1953 51 -1887 85
rect -1953 17 -1937 51
rect -1903 17 -1887 51
rect -1953 -17 -1887 17
rect -1953 -51 -1937 -17
rect -1903 -51 -1887 -17
rect -1953 -85 -1887 -51
rect -1953 -119 -1937 -85
rect -1903 -119 -1887 -85
rect -1953 -153 -1887 -119
rect -1953 -187 -1937 -153
rect -1903 -187 -1887 -153
rect -1953 -221 -1887 -187
rect -1953 -255 -1937 -221
rect -1903 -255 -1887 -221
rect -1953 -300 -1887 -255
rect -1857 255 -1791 300
rect -1857 221 -1841 255
rect -1807 221 -1791 255
rect -1857 187 -1791 221
rect -1857 153 -1841 187
rect -1807 153 -1791 187
rect -1857 119 -1791 153
rect -1857 85 -1841 119
rect -1807 85 -1791 119
rect -1857 51 -1791 85
rect -1857 17 -1841 51
rect -1807 17 -1791 51
rect -1857 -17 -1791 17
rect -1857 -51 -1841 -17
rect -1807 -51 -1791 -17
rect -1857 -85 -1791 -51
rect -1857 -119 -1841 -85
rect -1807 -119 -1791 -85
rect -1857 -153 -1791 -119
rect -1857 -187 -1841 -153
rect -1807 -187 -1791 -153
rect -1857 -221 -1791 -187
rect -1857 -255 -1841 -221
rect -1807 -255 -1791 -221
rect -1857 -300 -1791 -255
rect -1761 255 -1695 300
rect -1761 221 -1745 255
rect -1711 221 -1695 255
rect -1761 187 -1695 221
rect -1761 153 -1745 187
rect -1711 153 -1695 187
rect -1761 119 -1695 153
rect -1761 85 -1745 119
rect -1711 85 -1695 119
rect -1761 51 -1695 85
rect -1761 17 -1745 51
rect -1711 17 -1695 51
rect -1761 -17 -1695 17
rect -1761 -51 -1745 -17
rect -1711 -51 -1695 -17
rect -1761 -85 -1695 -51
rect -1761 -119 -1745 -85
rect -1711 -119 -1695 -85
rect -1761 -153 -1695 -119
rect -1761 -187 -1745 -153
rect -1711 -187 -1695 -153
rect -1761 -221 -1695 -187
rect -1761 -255 -1745 -221
rect -1711 -255 -1695 -221
rect -1761 -300 -1695 -255
rect -1665 255 -1599 300
rect -1665 221 -1649 255
rect -1615 221 -1599 255
rect -1665 187 -1599 221
rect -1665 153 -1649 187
rect -1615 153 -1599 187
rect -1665 119 -1599 153
rect -1665 85 -1649 119
rect -1615 85 -1599 119
rect -1665 51 -1599 85
rect -1665 17 -1649 51
rect -1615 17 -1599 51
rect -1665 -17 -1599 17
rect -1665 -51 -1649 -17
rect -1615 -51 -1599 -17
rect -1665 -85 -1599 -51
rect -1665 -119 -1649 -85
rect -1615 -119 -1599 -85
rect -1665 -153 -1599 -119
rect -1665 -187 -1649 -153
rect -1615 -187 -1599 -153
rect -1665 -221 -1599 -187
rect -1665 -255 -1649 -221
rect -1615 -255 -1599 -221
rect -1665 -300 -1599 -255
rect -1569 255 -1503 300
rect -1569 221 -1553 255
rect -1519 221 -1503 255
rect -1569 187 -1503 221
rect -1569 153 -1553 187
rect -1519 153 -1503 187
rect -1569 119 -1503 153
rect -1569 85 -1553 119
rect -1519 85 -1503 119
rect -1569 51 -1503 85
rect -1569 17 -1553 51
rect -1519 17 -1503 51
rect -1569 -17 -1503 17
rect -1569 -51 -1553 -17
rect -1519 -51 -1503 -17
rect -1569 -85 -1503 -51
rect -1569 -119 -1553 -85
rect -1519 -119 -1503 -85
rect -1569 -153 -1503 -119
rect -1569 -187 -1553 -153
rect -1519 -187 -1503 -153
rect -1569 -221 -1503 -187
rect -1569 -255 -1553 -221
rect -1519 -255 -1503 -221
rect -1569 -300 -1503 -255
rect -1473 255 -1407 300
rect -1473 221 -1457 255
rect -1423 221 -1407 255
rect -1473 187 -1407 221
rect -1473 153 -1457 187
rect -1423 153 -1407 187
rect -1473 119 -1407 153
rect -1473 85 -1457 119
rect -1423 85 -1407 119
rect -1473 51 -1407 85
rect -1473 17 -1457 51
rect -1423 17 -1407 51
rect -1473 -17 -1407 17
rect -1473 -51 -1457 -17
rect -1423 -51 -1407 -17
rect -1473 -85 -1407 -51
rect -1473 -119 -1457 -85
rect -1423 -119 -1407 -85
rect -1473 -153 -1407 -119
rect -1473 -187 -1457 -153
rect -1423 -187 -1407 -153
rect -1473 -221 -1407 -187
rect -1473 -255 -1457 -221
rect -1423 -255 -1407 -221
rect -1473 -300 -1407 -255
rect -1377 255 -1311 300
rect -1377 221 -1361 255
rect -1327 221 -1311 255
rect -1377 187 -1311 221
rect -1377 153 -1361 187
rect -1327 153 -1311 187
rect -1377 119 -1311 153
rect -1377 85 -1361 119
rect -1327 85 -1311 119
rect -1377 51 -1311 85
rect -1377 17 -1361 51
rect -1327 17 -1311 51
rect -1377 -17 -1311 17
rect -1377 -51 -1361 -17
rect -1327 -51 -1311 -17
rect -1377 -85 -1311 -51
rect -1377 -119 -1361 -85
rect -1327 -119 -1311 -85
rect -1377 -153 -1311 -119
rect -1377 -187 -1361 -153
rect -1327 -187 -1311 -153
rect -1377 -221 -1311 -187
rect -1377 -255 -1361 -221
rect -1327 -255 -1311 -221
rect -1377 -300 -1311 -255
rect -1281 255 -1215 300
rect -1281 221 -1265 255
rect -1231 221 -1215 255
rect -1281 187 -1215 221
rect -1281 153 -1265 187
rect -1231 153 -1215 187
rect -1281 119 -1215 153
rect -1281 85 -1265 119
rect -1231 85 -1215 119
rect -1281 51 -1215 85
rect -1281 17 -1265 51
rect -1231 17 -1215 51
rect -1281 -17 -1215 17
rect -1281 -51 -1265 -17
rect -1231 -51 -1215 -17
rect -1281 -85 -1215 -51
rect -1281 -119 -1265 -85
rect -1231 -119 -1215 -85
rect -1281 -153 -1215 -119
rect -1281 -187 -1265 -153
rect -1231 -187 -1215 -153
rect -1281 -221 -1215 -187
rect -1281 -255 -1265 -221
rect -1231 -255 -1215 -221
rect -1281 -300 -1215 -255
rect -1185 255 -1119 300
rect -1185 221 -1169 255
rect -1135 221 -1119 255
rect -1185 187 -1119 221
rect -1185 153 -1169 187
rect -1135 153 -1119 187
rect -1185 119 -1119 153
rect -1185 85 -1169 119
rect -1135 85 -1119 119
rect -1185 51 -1119 85
rect -1185 17 -1169 51
rect -1135 17 -1119 51
rect -1185 -17 -1119 17
rect -1185 -51 -1169 -17
rect -1135 -51 -1119 -17
rect -1185 -85 -1119 -51
rect -1185 -119 -1169 -85
rect -1135 -119 -1119 -85
rect -1185 -153 -1119 -119
rect -1185 -187 -1169 -153
rect -1135 -187 -1119 -153
rect -1185 -221 -1119 -187
rect -1185 -255 -1169 -221
rect -1135 -255 -1119 -221
rect -1185 -300 -1119 -255
rect -1089 255 -1023 300
rect -1089 221 -1073 255
rect -1039 221 -1023 255
rect -1089 187 -1023 221
rect -1089 153 -1073 187
rect -1039 153 -1023 187
rect -1089 119 -1023 153
rect -1089 85 -1073 119
rect -1039 85 -1023 119
rect -1089 51 -1023 85
rect -1089 17 -1073 51
rect -1039 17 -1023 51
rect -1089 -17 -1023 17
rect -1089 -51 -1073 -17
rect -1039 -51 -1023 -17
rect -1089 -85 -1023 -51
rect -1089 -119 -1073 -85
rect -1039 -119 -1023 -85
rect -1089 -153 -1023 -119
rect -1089 -187 -1073 -153
rect -1039 -187 -1023 -153
rect -1089 -221 -1023 -187
rect -1089 -255 -1073 -221
rect -1039 -255 -1023 -221
rect -1089 -300 -1023 -255
rect -993 255 -927 300
rect -993 221 -977 255
rect -943 221 -927 255
rect -993 187 -927 221
rect -993 153 -977 187
rect -943 153 -927 187
rect -993 119 -927 153
rect -993 85 -977 119
rect -943 85 -927 119
rect -993 51 -927 85
rect -993 17 -977 51
rect -943 17 -927 51
rect -993 -17 -927 17
rect -993 -51 -977 -17
rect -943 -51 -927 -17
rect -993 -85 -927 -51
rect -993 -119 -977 -85
rect -943 -119 -927 -85
rect -993 -153 -927 -119
rect -993 -187 -977 -153
rect -943 -187 -927 -153
rect -993 -221 -927 -187
rect -993 -255 -977 -221
rect -943 -255 -927 -221
rect -993 -300 -927 -255
rect -897 255 -831 300
rect -897 221 -881 255
rect -847 221 -831 255
rect -897 187 -831 221
rect -897 153 -881 187
rect -847 153 -831 187
rect -897 119 -831 153
rect -897 85 -881 119
rect -847 85 -831 119
rect -897 51 -831 85
rect -897 17 -881 51
rect -847 17 -831 51
rect -897 -17 -831 17
rect -897 -51 -881 -17
rect -847 -51 -831 -17
rect -897 -85 -831 -51
rect -897 -119 -881 -85
rect -847 -119 -831 -85
rect -897 -153 -831 -119
rect -897 -187 -881 -153
rect -847 -187 -831 -153
rect -897 -221 -831 -187
rect -897 -255 -881 -221
rect -847 -255 -831 -221
rect -897 -300 -831 -255
rect -801 255 -735 300
rect -801 221 -785 255
rect -751 221 -735 255
rect -801 187 -735 221
rect -801 153 -785 187
rect -751 153 -735 187
rect -801 119 -735 153
rect -801 85 -785 119
rect -751 85 -735 119
rect -801 51 -735 85
rect -801 17 -785 51
rect -751 17 -735 51
rect -801 -17 -735 17
rect -801 -51 -785 -17
rect -751 -51 -735 -17
rect -801 -85 -735 -51
rect -801 -119 -785 -85
rect -751 -119 -735 -85
rect -801 -153 -735 -119
rect -801 -187 -785 -153
rect -751 -187 -735 -153
rect -801 -221 -735 -187
rect -801 -255 -785 -221
rect -751 -255 -735 -221
rect -801 -300 -735 -255
rect -705 255 -639 300
rect -705 221 -689 255
rect -655 221 -639 255
rect -705 187 -639 221
rect -705 153 -689 187
rect -655 153 -639 187
rect -705 119 -639 153
rect -705 85 -689 119
rect -655 85 -639 119
rect -705 51 -639 85
rect -705 17 -689 51
rect -655 17 -639 51
rect -705 -17 -639 17
rect -705 -51 -689 -17
rect -655 -51 -639 -17
rect -705 -85 -639 -51
rect -705 -119 -689 -85
rect -655 -119 -639 -85
rect -705 -153 -639 -119
rect -705 -187 -689 -153
rect -655 -187 -639 -153
rect -705 -221 -639 -187
rect -705 -255 -689 -221
rect -655 -255 -639 -221
rect -705 -300 -639 -255
rect -609 255 -543 300
rect -609 221 -593 255
rect -559 221 -543 255
rect -609 187 -543 221
rect -609 153 -593 187
rect -559 153 -543 187
rect -609 119 -543 153
rect -609 85 -593 119
rect -559 85 -543 119
rect -609 51 -543 85
rect -609 17 -593 51
rect -559 17 -543 51
rect -609 -17 -543 17
rect -609 -51 -593 -17
rect -559 -51 -543 -17
rect -609 -85 -543 -51
rect -609 -119 -593 -85
rect -559 -119 -543 -85
rect -609 -153 -543 -119
rect -609 -187 -593 -153
rect -559 -187 -543 -153
rect -609 -221 -543 -187
rect -609 -255 -593 -221
rect -559 -255 -543 -221
rect -609 -300 -543 -255
rect -513 255 -447 300
rect -513 221 -497 255
rect -463 221 -447 255
rect -513 187 -447 221
rect -513 153 -497 187
rect -463 153 -447 187
rect -513 119 -447 153
rect -513 85 -497 119
rect -463 85 -447 119
rect -513 51 -447 85
rect -513 17 -497 51
rect -463 17 -447 51
rect -513 -17 -447 17
rect -513 -51 -497 -17
rect -463 -51 -447 -17
rect -513 -85 -447 -51
rect -513 -119 -497 -85
rect -463 -119 -447 -85
rect -513 -153 -447 -119
rect -513 -187 -497 -153
rect -463 -187 -447 -153
rect -513 -221 -447 -187
rect -513 -255 -497 -221
rect -463 -255 -447 -221
rect -513 -300 -447 -255
rect -417 255 -351 300
rect -417 221 -401 255
rect -367 221 -351 255
rect -417 187 -351 221
rect -417 153 -401 187
rect -367 153 -351 187
rect -417 119 -351 153
rect -417 85 -401 119
rect -367 85 -351 119
rect -417 51 -351 85
rect -417 17 -401 51
rect -367 17 -351 51
rect -417 -17 -351 17
rect -417 -51 -401 -17
rect -367 -51 -351 -17
rect -417 -85 -351 -51
rect -417 -119 -401 -85
rect -367 -119 -351 -85
rect -417 -153 -351 -119
rect -417 -187 -401 -153
rect -367 -187 -351 -153
rect -417 -221 -351 -187
rect -417 -255 -401 -221
rect -367 -255 -351 -221
rect -417 -300 -351 -255
rect -321 255 -255 300
rect -321 221 -305 255
rect -271 221 -255 255
rect -321 187 -255 221
rect -321 153 -305 187
rect -271 153 -255 187
rect -321 119 -255 153
rect -321 85 -305 119
rect -271 85 -255 119
rect -321 51 -255 85
rect -321 17 -305 51
rect -271 17 -255 51
rect -321 -17 -255 17
rect -321 -51 -305 -17
rect -271 -51 -255 -17
rect -321 -85 -255 -51
rect -321 -119 -305 -85
rect -271 -119 -255 -85
rect -321 -153 -255 -119
rect -321 -187 -305 -153
rect -271 -187 -255 -153
rect -321 -221 -255 -187
rect -321 -255 -305 -221
rect -271 -255 -255 -221
rect -321 -300 -255 -255
rect -225 255 -159 300
rect -225 221 -209 255
rect -175 221 -159 255
rect -225 187 -159 221
rect -225 153 -209 187
rect -175 153 -159 187
rect -225 119 -159 153
rect -225 85 -209 119
rect -175 85 -159 119
rect -225 51 -159 85
rect -225 17 -209 51
rect -175 17 -159 51
rect -225 -17 -159 17
rect -225 -51 -209 -17
rect -175 -51 -159 -17
rect -225 -85 -159 -51
rect -225 -119 -209 -85
rect -175 -119 -159 -85
rect -225 -153 -159 -119
rect -225 -187 -209 -153
rect -175 -187 -159 -153
rect -225 -221 -159 -187
rect -225 -255 -209 -221
rect -175 -255 -159 -221
rect -225 -300 -159 -255
rect -129 255 -63 300
rect -129 221 -113 255
rect -79 221 -63 255
rect -129 187 -63 221
rect -129 153 -113 187
rect -79 153 -63 187
rect -129 119 -63 153
rect -129 85 -113 119
rect -79 85 -63 119
rect -129 51 -63 85
rect -129 17 -113 51
rect -79 17 -63 51
rect -129 -17 -63 17
rect -129 -51 -113 -17
rect -79 -51 -63 -17
rect -129 -85 -63 -51
rect -129 -119 -113 -85
rect -79 -119 -63 -85
rect -129 -153 -63 -119
rect -129 -187 -113 -153
rect -79 -187 -63 -153
rect -129 -221 -63 -187
rect -129 -255 -113 -221
rect -79 -255 -63 -221
rect -129 -300 -63 -255
rect -33 255 33 300
rect -33 221 -17 255
rect 17 221 33 255
rect -33 187 33 221
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -221 33 -187
rect -33 -255 -17 -221
rect 17 -255 33 -221
rect -33 -300 33 -255
rect 63 255 129 300
rect 63 221 79 255
rect 113 221 129 255
rect 63 187 129 221
rect 63 153 79 187
rect 113 153 129 187
rect 63 119 129 153
rect 63 85 79 119
rect 113 85 129 119
rect 63 51 129 85
rect 63 17 79 51
rect 113 17 129 51
rect 63 -17 129 17
rect 63 -51 79 -17
rect 113 -51 129 -17
rect 63 -85 129 -51
rect 63 -119 79 -85
rect 113 -119 129 -85
rect 63 -153 129 -119
rect 63 -187 79 -153
rect 113 -187 129 -153
rect 63 -221 129 -187
rect 63 -255 79 -221
rect 113 -255 129 -221
rect 63 -300 129 -255
rect 159 255 225 300
rect 159 221 175 255
rect 209 221 225 255
rect 159 187 225 221
rect 159 153 175 187
rect 209 153 225 187
rect 159 119 225 153
rect 159 85 175 119
rect 209 85 225 119
rect 159 51 225 85
rect 159 17 175 51
rect 209 17 225 51
rect 159 -17 225 17
rect 159 -51 175 -17
rect 209 -51 225 -17
rect 159 -85 225 -51
rect 159 -119 175 -85
rect 209 -119 225 -85
rect 159 -153 225 -119
rect 159 -187 175 -153
rect 209 -187 225 -153
rect 159 -221 225 -187
rect 159 -255 175 -221
rect 209 -255 225 -221
rect 159 -300 225 -255
rect 255 255 321 300
rect 255 221 271 255
rect 305 221 321 255
rect 255 187 321 221
rect 255 153 271 187
rect 305 153 321 187
rect 255 119 321 153
rect 255 85 271 119
rect 305 85 321 119
rect 255 51 321 85
rect 255 17 271 51
rect 305 17 321 51
rect 255 -17 321 17
rect 255 -51 271 -17
rect 305 -51 321 -17
rect 255 -85 321 -51
rect 255 -119 271 -85
rect 305 -119 321 -85
rect 255 -153 321 -119
rect 255 -187 271 -153
rect 305 -187 321 -153
rect 255 -221 321 -187
rect 255 -255 271 -221
rect 305 -255 321 -221
rect 255 -300 321 -255
rect 351 255 417 300
rect 351 221 367 255
rect 401 221 417 255
rect 351 187 417 221
rect 351 153 367 187
rect 401 153 417 187
rect 351 119 417 153
rect 351 85 367 119
rect 401 85 417 119
rect 351 51 417 85
rect 351 17 367 51
rect 401 17 417 51
rect 351 -17 417 17
rect 351 -51 367 -17
rect 401 -51 417 -17
rect 351 -85 417 -51
rect 351 -119 367 -85
rect 401 -119 417 -85
rect 351 -153 417 -119
rect 351 -187 367 -153
rect 401 -187 417 -153
rect 351 -221 417 -187
rect 351 -255 367 -221
rect 401 -255 417 -221
rect 351 -300 417 -255
rect 447 255 513 300
rect 447 221 463 255
rect 497 221 513 255
rect 447 187 513 221
rect 447 153 463 187
rect 497 153 513 187
rect 447 119 513 153
rect 447 85 463 119
rect 497 85 513 119
rect 447 51 513 85
rect 447 17 463 51
rect 497 17 513 51
rect 447 -17 513 17
rect 447 -51 463 -17
rect 497 -51 513 -17
rect 447 -85 513 -51
rect 447 -119 463 -85
rect 497 -119 513 -85
rect 447 -153 513 -119
rect 447 -187 463 -153
rect 497 -187 513 -153
rect 447 -221 513 -187
rect 447 -255 463 -221
rect 497 -255 513 -221
rect 447 -300 513 -255
rect 543 255 609 300
rect 543 221 559 255
rect 593 221 609 255
rect 543 187 609 221
rect 543 153 559 187
rect 593 153 609 187
rect 543 119 609 153
rect 543 85 559 119
rect 593 85 609 119
rect 543 51 609 85
rect 543 17 559 51
rect 593 17 609 51
rect 543 -17 609 17
rect 543 -51 559 -17
rect 593 -51 609 -17
rect 543 -85 609 -51
rect 543 -119 559 -85
rect 593 -119 609 -85
rect 543 -153 609 -119
rect 543 -187 559 -153
rect 593 -187 609 -153
rect 543 -221 609 -187
rect 543 -255 559 -221
rect 593 -255 609 -221
rect 543 -300 609 -255
rect 639 255 705 300
rect 639 221 655 255
rect 689 221 705 255
rect 639 187 705 221
rect 639 153 655 187
rect 689 153 705 187
rect 639 119 705 153
rect 639 85 655 119
rect 689 85 705 119
rect 639 51 705 85
rect 639 17 655 51
rect 689 17 705 51
rect 639 -17 705 17
rect 639 -51 655 -17
rect 689 -51 705 -17
rect 639 -85 705 -51
rect 639 -119 655 -85
rect 689 -119 705 -85
rect 639 -153 705 -119
rect 639 -187 655 -153
rect 689 -187 705 -153
rect 639 -221 705 -187
rect 639 -255 655 -221
rect 689 -255 705 -221
rect 639 -300 705 -255
rect 735 255 801 300
rect 735 221 751 255
rect 785 221 801 255
rect 735 187 801 221
rect 735 153 751 187
rect 785 153 801 187
rect 735 119 801 153
rect 735 85 751 119
rect 785 85 801 119
rect 735 51 801 85
rect 735 17 751 51
rect 785 17 801 51
rect 735 -17 801 17
rect 735 -51 751 -17
rect 785 -51 801 -17
rect 735 -85 801 -51
rect 735 -119 751 -85
rect 785 -119 801 -85
rect 735 -153 801 -119
rect 735 -187 751 -153
rect 785 -187 801 -153
rect 735 -221 801 -187
rect 735 -255 751 -221
rect 785 -255 801 -221
rect 735 -300 801 -255
rect 831 255 897 300
rect 831 221 847 255
rect 881 221 897 255
rect 831 187 897 221
rect 831 153 847 187
rect 881 153 897 187
rect 831 119 897 153
rect 831 85 847 119
rect 881 85 897 119
rect 831 51 897 85
rect 831 17 847 51
rect 881 17 897 51
rect 831 -17 897 17
rect 831 -51 847 -17
rect 881 -51 897 -17
rect 831 -85 897 -51
rect 831 -119 847 -85
rect 881 -119 897 -85
rect 831 -153 897 -119
rect 831 -187 847 -153
rect 881 -187 897 -153
rect 831 -221 897 -187
rect 831 -255 847 -221
rect 881 -255 897 -221
rect 831 -300 897 -255
rect 927 255 993 300
rect 927 221 943 255
rect 977 221 993 255
rect 927 187 993 221
rect 927 153 943 187
rect 977 153 993 187
rect 927 119 993 153
rect 927 85 943 119
rect 977 85 993 119
rect 927 51 993 85
rect 927 17 943 51
rect 977 17 993 51
rect 927 -17 993 17
rect 927 -51 943 -17
rect 977 -51 993 -17
rect 927 -85 993 -51
rect 927 -119 943 -85
rect 977 -119 993 -85
rect 927 -153 993 -119
rect 927 -187 943 -153
rect 977 -187 993 -153
rect 927 -221 993 -187
rect 927 -255 943 -221
rect 977 -255 993 -221
rect 927 -300 993 -255
rect 1023 255 1089 300
rect 1023 221 1039 255
rect 1073 221 1089 255
rect 1023 187 1089 221
rect 1023 153 1039 187
rect 1073 153 1089 187
rect 1023 119 1089 153
rect 1023 85 1039 119
rect 1073 85 1089 119
rect 1023 51 1089 85
rect 1023 17 1039 51
rect 1073 17 1089 51
rect 1023 -17 1089 17
rect 1023 -51 1039 -17
rect 1073 -51 1089 -17
rect 1023 -85 1089 -51
rect 1023 -119 1039 -85
rect 1073 -119 1089 -85
rect 1023 -153 1089 -119
rect 1023 -187 1039 -153
rect 1073 -187 1089 -153
rect 1023 -221 1089 -187
rect 1023 -255 1039 -221
rect 1073 -255 1089 -221
rect 1023 -300 1089 -255
rect 1119 255 1185 300
rect 1119 221 1135 255
rect 1169 221 1185 255
rect 1119 187 1185 221
rect 1119 153 1135 187
rect 1169 153 1185 187
rect 1119 119 1185 153
rect 1119 85 1135 119
rect 1169 85 1185 119
rect 1119 51 1185 85
rect 1119 17 1135 51
rect 1169 17 1185 51
rect 1119 -17 1185 17
rect 1119 -51 1135 -17
rect 1169 -51 1185 -17
rect 1119 -85 1185 -51
rect 1119 -119 1135 -85
rect 1169 -119 1185 -85
rect 1119 -153 1185 -119
rect 1119 -187 1135 -153
rect 1169 -187 1185 -153
rect 1119 -221 1185 -187
rect 1119 -255 1135 -221
rect 1169 -255 1185 -221
rect 1119 -300 1185 -255
rect 1215 255 1281 300
rect 1215 221 1231 255
rect 1265 221 1281 255
rect 1215 187 1281 221
rect 1215 153 1231 187
rect 1265 153 1281 187
rect 1215 119 1281 153
rect 1215 85 1231 119
rect 1265 85 1281 119
rect 1215 51 1281 85
rect 1215 17 1231 51
rect 1265 17 1281 51
rect 1215 -17 1281 17
rect 1215 -51 1231 -17
rect 1265 -51 1281 -17
rect 1215 -85 1281 -51
rect 1215 -119 1231 -85
rect 1265 -119 1281 -85
rect 1215 -153 1281 -119
rect 1215 -187 1231 -153
rect 1265 -187 1281 -153
rect 1215 -221 1281 -187
rect 1215 -255 1231 -221
rect 1265 -255 1281 -221
rect 1215 -300 1281 -255
rect 1311 255 1377 300
rect 1311 221 1327 255
rect 1361 221 1377 255
rect 1311 187 1377 221
rect 1311 153 1327 187
rect 1361 153 1377 187
rect 1311 119 1377 153
rect 1311 85 1327 119
rect 1361 85 1377 119
rect 1311 51 1377 85
rect 1311 17 1327 51
rect 1361 17 1377 51
rect 1311 -17 1377 17
rect 1311 -51 1327 -17
rect 1361 -51 1377 -17
rect 1311 -85 1377 -51
rect 1311 -119 1327 -85
rect 1361 -119 1377 -85
rect 1311 -153 1377 -119
rect 1311 -187 1327 -153
rect 1361 -187 1377 -153
rect 1311 -221 1377 -187
rect 1311 -255 1327 -221
rect 1361 -255 1377 -221
rect 1311 -300 1377 -255
rect 1407 255 1473 300
rect 1407 221 1423 255
rect 1457 221 1473 255
rect 1407 187 1473 221
rect 1407 153 1423 187
rect 1457 153 1473 187
rect 1407 119 1473 153
rect 1407 85 1423 119
rect 1457 85 1473 119
rect 1407 51 1473 85
rect 1407 17 1423 51
rect 1457 17 1473 51
rect 1407 -17 1473 17
rect 1407 -51 1423 -17
rect 1457 -51 1473 -17
rect 1407 -85 1473 -51
rect 1407 -119 1423 -85
rect 1457 -119 1473 -85
rect 1407 -153 1473 -119
rect 1407 -187 1423 -153
rect 1457 -187 1473 -153
rect 1407 -221 1473 -187
rect 1407 -255 1423 -221
rect 1457 -255 1473 -221
rect 1407 -300 1473 -255
rect 1503 255 1569 300
rect 1503 221 1519 255
rect 1553 221 1569 255
rect 1503 187 1569 221
rect 1503 153 1519 187
rect 1553 153 1569 187
rect 1503 119 1569 153
rect 1503 85 1519 119
rect 1553 85 1569 119
rect 1503 51 1569 85
rect 1503 17 1519 51
rect 1553 17 1569 51
rect 1503 -17 1569 17
rect 1503 -51 1519 -17
rect 1553 -51 1569 -17
rect 1503 -85 1569 -51
rect 1503 -119 1519 -85
rect 1553 -119 1569 -85
rect 1503 -153 1569 -119
rect 1503 -187 1519 -153
rect 1553 -187 1569 -153
rect 1503 -221 1569 -187
rect 1503 -255 1519 -221
rect 1553 -255 1569 -221
rect 1503 -300 1569 -255
rect 1599 255 1665 300
rect 1599 221 1615 255
rect 1649 221 1665 255
rect 1599 187 1665 221
rect 1599 153 1615 187
rect 1649 153 1665 187
rect 1599 119 1665 153
rect 1599 85 1615 119
rect 1649 85 1665 119
rect 1599 51 1665 85
rect 1599 17 1615 51
rect 1649 17 1665 51
rect 1599 -17 1665 17
rect 1599 -51 1615 -17
rect 1649 -51 1665 -17
rect 1599 -85 1665 -51
rect 1599 -119 1615 -85
rect 1649 -119 1665 -85
rect 1599 -153 1665 -119
rect 1599 -187 1615 -153
rect 1649 -187 1665 -153
rect 1599 -221 1665 -187
rect 1599 -255 1615 -221
rect 1649 -255 1665 -221
rect 1599 -300 1665 -255
rect 1695 255 1761 300
rect 1695 221 1711 255
rect 1745 221 1761 255
rect 1695 187 1761 221
rect 1695 153 1711 187
rect 1745 153 1761 187
rect 1695 119 1761 153
rect 1695 85 1711 119
rect 1745 85 1761 119
rect 1695 51 1761 85
rect 1695 17 1711 51
rect 1745 17 1761 51
rect 1695 -17 1761 17
rect 1695 -51 1711 -17
rect 1745 -51 1761 -17
rect 1695 -85 1761 -51
rect 1695 -119 1711 -85
rect 1745 -119 1761 -85
rect 1695 -153 1761 -119
rect 1695 -187 1711 -153
rect 1745 -187 1761 -153
rect 1695 -221 1761 -187
rect 1695 -255 1711 -221
rect 1745 -255 1761 -221
rect 1695 -300 1761 -255
rect 1791 255 1857 300
rect 1791 221 1807 255
rect 1841 221 1857 255
rect 1791 187 1857 221
rect 1791 153 1807 187
rect 1841 153 1857 187
rect 1791 119 1857 153
rect 1791 85 1807 119
rect 1841 85 1857 119
rect 1791 51 1857 85
rect 1791 17 1807 51
rect 1841 17 1857 51
rect 1791 -17 1857 17
rect 1791 -51 1807 -17
rect 1841 -51 1857 -17
rect 1791 -85 1857 -51
rect 1791 -119 1807 -85
rect 1841 -119 1857 -85
rect 1791 -153 1857 -119
rect 1791 -187 1807 -153
rect 1841 -187 1857 -153
rect 1791 -221 1857 -187
rect 1791 -255 1807 -221
rect 1841 -255 1857 -221
rect 1791 -300 1857 -255
rect 1887 255 1953 300
rect 1887 221 1903 255
rect 1937 221 1953 255
rect 1887 187 1953 221
rect 1887 153 1903 187
rect 1937 153 1953 187
rect 1887 119 1953 153
rect 1887 85 1903 119
rect 1937 85 1953 119
rect 1887 51 1953 85
rect 1887 17 1903 51
rect 1937 17 1953 51
rect 1887 -17 1953 17
rect 1887 -51 1903 -17
rect 1937 -51 1953 -17
rect 1887 -85 1953 -51
rect 1887 -119 1903 -85
rect 1937 -119 1953 -85
rect 1887 -153 1953 -119
rect 1887 -187 1903 -153
rect 1937 -187 1953 -153
rect 1887 -221 1953 -187
rect 1887 -255 1903 -221
rect 1937 -255 1953 -221
rect 1887 -300 1953 -255
rect 1983 255 2045 300
rect 1983 221 1999 255
rect 2033 221 2045 255
rect 1983 187 2045 221
rect 1983 153 1999 187
rect 2033 153 2045 187
rect 1983 119 2045 153
rect 1983 85 1999 119
rect 2033 85 2045 119
rect 1983 51 2045 85
rect 1983 17 1999 51
rect 2033 17 2045 51
rect 1983 -17 2045 17
rect 1983 -51 1999 -17
rect 2033 -51 2045 -17
rect 1983 -85 2045 -51
rect 1983 -119 1999 -85
rect 2033 -119 2045 -85
rect 1983 -153 2045 -119
rect 1983 -187 1999 -153
rect 2033 -187 2045 -153
rect 1983 -221 2045 -187
rect 1983 -255 1999 -221
rect 2033 -255 2045 -221
rect 1983 -300 2045 -255
<< pdiffc >>
rect -2033 221 -1999 255
rect -2033 153 -1999 187
rect -2033 85 -1999 119
rect -2033 17 -1999 51
rect -2033 -51 -1999 -17
rect -2033 -119 -1999 -85
rect -2033 -187 -1999 -153
rect -2033 -255 -1999 -221
rect -1937 221 -1903 255
rect -1937 153 -1903 187
rect -1937 85 -1903 119
rect -1937 17 -1903 51
rect -1937 -51 -1903 -17
rect -1937 -119 -1903 -85
rect -1937 -187 -1903 -153
rect -1937 -255 -1903 -221
rect -1841 221 -1807 255
rect -1841 153 -1807 187
rect -1841 85 -1807 119
rect -1841 17 -1807 51
rect -1841 -51 -1807 -17
rect -1841 -119 -1807 -85
rect -1841 -187 -1807 -153
rect -1841 -255 -1807 -221
rect -1745 221 -1711 255
rect -1745 153 -1711 187
rect -1745 85 -1711 119
rect -1745 17 -1711 51
rect -1745 -51 -1711 -17
rect -1745 -119 -1711 -85
rect -1745 -187 -1711 -153
rect -1745 -255 -1711 -221
rect -1649 221 -1615 255
rect -1649 153 -1615 187
rect -1649 85 -1615 119
rect -1649 17 -1615 51
rect -1649 -51 -1615 -17
rect -1649 -119 -1615 -85
rect -1649 -187 -1615 -153
rect -1649 -255 -1615 -221
rect -1553 221 -1519 255
rect -1553 153 -1519 187
rect -1553 85 -1519 119
rect -1553 17 -1519 51
rect -1553 -51 -1519 -17
rect -1553 -119 -1519 -85
rect -1553 -187 -1519 -153
rect -1553 -255 -1519 -221
rect -1457 221 -1423 255
rect -1457 153 -1423 187
rect -1457 85 -1423 119
rect -1457 17 -1423 51
rect -1457 -51 -1423 -17
rect -1457 -119 -1423 -85
rect -1457 -187 -1423 -153
rect -1457 -255 -1423 -221
rect -1361 221 -1327 255
rect -1361 153 -1327 187
rect -1361 85 -1327 119
rect -1361 17 -1327 51
rect -1361 -51 -1327 -17
rect -1361 -119 -1327 -85
rect -1361 -187 -1327 -153
rect -1361 -255 -1327 -221
rect -1265 221 -1231 255
rect -1265 153 -1231 187
rect -1265 85 -1231 119
rect -1265 17 -1231 51
rect -1265 -51 -1231 -17
rect -1265 -119 -1231 -85
rect -1265 -187 -1231 -153
rect -1265 -255 -1231 -221
rect -1169 221 -1135 255
rect -1169 153 -1135 187
rect -1169 85 -1135 119
rect -1169 17 -1135 51
rect -1169 -51 -1135 -17
rect -1169 -119 -1135 -85
rect -1169 -187 -1135 -153
rect -1169 -255 -1135 -221
rect -1073 221 -1039 255
rect -1073 153 -1039 187
rect -1073 85 -1039 119
rect -1073 17 -1039 51
rect -1073 -51 -1039 -17
rect -1073 -119 -1039 -85
rect -1073 -187 -1039 -153
rect -1073 -255 -1039 -221
rect -977 221 -943 255
rect -977 153 -943 187
rect -977 85 -943 119
rect -977 17 -943 51
rect -977 -51 -943 -17
rect -977 -119 -943 -85
rect -977 -187 -943 -153
rect -977 -255 -943 -221
rect -881 221 -847 255
rect -881 153 -847 187
rect -881 85 -847 119
rect -881 17 -847 51
rect -881 -51 -847 -17
rect -881 -119 -847 -85
rect -881 -187 -847 -153
rect -881 -255 -847 -221
rect -785 221 -751 255
rect -785 153 -751 187
rect -785 85 -751 119
rect -785 17 -751 51
rect -785 -51 -751 -17
rect -785 -119 -751 -85
rect -785 -187 -751 -153
rect -785 -255 -751 -221
rect -689 221 -655 255
rect -689 153 -655 187
rect -689 85 -655 119
rect -689 17 -655 51
rect -689 -51 -655 -17
rect -689 -119 -655 -85
rect -689 -187 -655 -153
rect -689 -255 -655 -221
rect -593 221 -559 255
rect -593 153 -559 187
rect -593 85 -559 119
rect -593 17 -559 51
rect -593 -51 -559 -17
rect -593 -119 -559 -85
rect -593 -187 -559 -153
rect -593 -255 -559 -221
rect -497 221 -463 255
rect -497 153 -463 187
rect -497 85 -463 119
rect -497 17 -463 51
rect -497 -51 -463 -17
rect -497 -119 -463 -85
rect -497 -187 -463 -153
rect -497 -255 -463 -221
rect -401 221 -367 255
rect -401 153 -367 187
rect -401 85 -367 119
rect -401 17 -367 51
rect -401 -51 -367 -17
rect -401 -119 -367 -85
rect -401 -187 -367 -153
rect -401 -255 -367 -221
rect -305 221 -271 255
rect -305 153 -271 187
rect -305 85 -271 119
rect -305 17 -271 51
rect -305 -51 -271 -17
rect -305 -119 -271 -85
rect -305 -187 -271 -153
rect -305 -255 -271 -221
rect -209 221 -175 255
rect -209 153 -175 187
rect -209 85 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -85
rect -209 -187 -175 -153
rect -209 -255 -175 -221
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 175 221 209 255
rect 175 153 209 187
rect 175 85 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -85
rect 175 -187 209 -153
rect 175 -255 209 -221
rect 271 221 305 255
rect 271 153 305 187
rect 271 85 305 119
rect 271 17 305 51
rect 271 -51 305 -17
rect 271 -119 305 -85
rect 271 -187 305 -153
rect 271 -255 305 -221
rect 367 221 401 255
rect 367 153 401 187
rect 367 85 401 119
rect 367 17 401 51
rect 367 -51 401 -17
rect 367 -119 401 -85
rect 367 -187 401 -153
rect 367 -255 401 -221
rect 463 221 497 255
rect 463 153 497 187
rect 463 85 497 119
rect 463 17 497 51
rect 463 -51 497 -17
rect 463 -119 497 -85
rect 463 -187 497 -153
rect 463 -255 497 -221
rect 559 221 593 255
rect 559 153 593 187
rect 559 85 593 119
rect 559 17 593 51
rect 559 -51 593 -17
rect 559 -119 593 -85
rect 559 -187 593 -153
rect 559 -255 593 -221
rect 655 221 689 255
rect 655 153 689 187
rect 655 85 689 119
rect 655 17 689 51
rect 655 -51 689 -17
rect 655 -119 689 -85
rect 655 -187 689 -153
rect 655 -255 689 -221
rect 751 221 785 255
rect 751 153 785 187
rect 751 85 785 119
rect 751 17 785 51
rect 751 -51 785 -17
rect 751 -119 785 -85
rect 751 -187 785 -153
rect 751 -255 785 -221
rect 847 221 881 255
rect 847 153 881 187
rect 847 85 881 119
rect 847 17 881 51
rect 847 -51 881 -17
rect 847 -119 881 -85
rect 847 -187 881 -153
rect 847 -255 881 -221
rect 943 221 977 255
rect 943 153 977 187
rect 943 85 977 119
rect 943 17 977 51
rect 943 -51 977 -17
rect 943 -119 977 -85
rect 943 -187 977 -153
rect 943 -255 977 -221
rect 1039 221 1073 255
rect 1039 153 1073 187
rect 1039 85 1073 119
rect 1039 17 1073 51
rect 1039 -51 1073 -17
rect 1039 -119 1073 -85
rect 1039 -187 1073 -153
rect 1039 -255 1073 -221
rect 1135 221 1169 255
rect 1135 153 1169 187
rect 1135 85 1169 119
rect 1135 17 1169 51
rect 1135 -51 1169 -17
rect 1135 -119 1169 -85
rect 1135 -187 1169 -153
rect 1135 -255 1169 -221
rect 1231 221 1265 255
rect 1231 153 1265 187
rect 1231 85 1265 119
rect 1231 17 1265 51
rect 1231 -51 1265 -17
rect 1231 -119 1265 -85
rect 1231 -187 1265 -153
rect 1231 -255 1265 -221
rect 1327 221 1361 255
rect 1327 153 1361 187
rect 1327 85 1361 119
rect 1327 17 1361 51
rect 1327 -51 1361 -17
rect 1327 -119 1361 -85
rect 1327 -187 1361 -153
rect 1327 -255 1361 -221
rect 1423 221 1457 255
rect 1423 153 1457 187
rect 1423 85 1457 119
rect 1423 17 1457 51
rect 1423 -51 1457 -17
rect 1423 -119 1457 -85
rect 1423 -187 1457 -153
rect 1423 -255 1457 -221
rect 1519 221 1553 255
rect 1519 153 1553 187
rect 1519 85 1553 119
rect 1519 17 1553 51
rect 1519 -51 1553 -17
rect 1519 -119 1553 -85
rect 1519 -187 1553 -153
rect 1519 -255 1553 -221
rect 1615 221 1649 255
rect 1615 153 1649 187
rect 1615 85 1649 119
rect 1615 17 1649 51
rect 1615 -51 1649 -17
rect 1615 -119 1649 -85
rect 1615 -187 1649 -153
rect 1615 -255 1649 -221
rect 1711 221 1745 255
rect 1711 153 1745 187
rect 1711 85 1745 119
rect 1711 17 1745 51
rect 1711 -51 1745 -17
rect 1711 -119 1745 -85
rect 1711 -187 1745 -153
rect 1711 -255 1745 -221
rect 1807 221 1841 255
rect 1807 153 1841 187
rect 1807 85 1841 119
rect 1807 17 1841 51
rect 1807 -51 1841 -17
rect 1807 -119 1841 -85
rect 1807 -187 1841 -153
rect 1807 -255 1841 -221
rect 1903 221 1937 255
rect 1903 153 1937 187
rect 1903 85 1937 119
rect 1903 17 1937 51
rect 1903 -51 1937 -17
rect 1903 -119 1937 -85
rect 1903 -187 1937 -153
rect 1903 -255 1937 -221
rect 1999 221 2033 255
rect 1999 153 2033 187
rect 1999 85 2033 119
rect 1999 17 2033 51
rect 1999 -51 2033 -17
rect 1999 -119 2033 -85
rect 1999 -187 2033 -153
rect 1999 -255 2033 -221
<< poly >>
rect -1905 381 -1839 397
rect -1905 347 -1889 381
rect -1855 347 -1839 381
rect -1905 331 -1839 347
rect -1713 381 -1647 397
rect -1713 347 -1697 381
rect -1663 347 -1647 381
rect -1713 331 -1647 347
rect -1521 381 -1455 397
rect -1521 347 -1505 381
rect -1471 347 -1455 381
rect -1521 331 -1455 347
rect -1329 381 -1263 397
rect -1329 347 -1313 381
rect -1279 347 -1263 381
rect -1329 331 -1263 347
rect -1137 381 -1071 397
rect -1137 347 -1121 381
rect -1087 347 -1071 381
rect -1137 331 -1071 347
rect -945 381 -879 397
rect -945 347 -929 381
rect -895 347 -879 381
rect -945 331 -879 347
rect -753 381 -687 397
rect -753 347 -737 381
rect -703 347 -687 381
rect -753 331 -687 347
rect -561 381 -495 397
rect -561 347 -545 381
rect -511 347 -495 381
rect -561 331 -495 347
rect -369 381 -303 397
rect -369 347 -353 381
rect -319 347 -303 381
rect -369 331 -303 347
rect -177 381 -111 397
rect -177 347 -161 381
rect -127 347 -111 381
rect -177 331 -111 347
rect 15 381 81 397
rect 15 347 31 381
rect 65 347 81 381
rect 15 331 81 347
rect 207 381 273 397
rect 207 347 223 381
rect 257 347 273 381
rect 207 331 273 347
rect 399 381 465 397
rect 399 347 415 381
rect 449 347 465 381
rect 399 331 465 347
rect 591 381 657 397
rect 591 347 607 381
rect 641 347 657 381
rect 591 331 657 347
rect 783 381 849 397
rect 783 347 799 381
rect 833 347 849 381
rect 783 331 849 347
rect 975 381 1041 397
rect 975 347 991 381
rect 1025 347 1041 381
rect 975 331 1041 347
rect 1167 381 1233 397
rect 1167 347 1183 381
rect 1217 347 1233 381
rect 1167 331 1233 347
rect 1359 381 1425 397
rect 1359 347 1375 381
rect 1409 347 1425 381
rect 1359 331 1425 347
rect 1551 381 1617 397
rect 1551 347 1567 381
rect 1601 347 1617 381
rect 1551 331 1617 347
rect 1743 381 1809 397
rect 1743 347 1759 381
rect 1793 347 1809 381
rect 1743 331 1809 347
rect 1935 381 2001 397
rect 1935 347 1951 381
rect 1985 347 2001 381
rect 1935 331 2001 347
rect -1983 300 -1953 326
rect -1887 300 -1857 331
rect -1791 300 -1761 326
rect -1695 300 -1665 331
rect -1599 300 -1569 326
rect -1503 300 -1473 331
rect -1407 300 -1377 326
rect -1311 300 -1281 331
rect -1215 300 -1185 326
rect -1119 300 -1089 331
rect -1023 300 -993 326
rect -927 300 -897 331
rect -831 300 -801 326
rect -735 300 -705 331
rect -639 300 -609 326
rect -543 300 -513 331
rect -447 300 -417 326
rect -351 300 -321 331
rect -255 300 -225 326
rect -159 300 -129 331
rect -63 300 -33 326
rect 33 300 63 331
rect 129 300 159 326
rect 225 300 255 331
rect 321 300 351 326
rect 417 300 447 331
rect 513 300 543 326
rect 609 300 639 331
rect 705 300 735 326
rect 801 300 831 331
rect 897 300 927 326
rect 993 300 1023 331
rect 1089 300 1119 326
rect 1185 300 1215 331
rect 1281 300 1311 326
rect 1377 300 1407 331
rect 1473 300 1503 326
rect 1569 300 1599 331
rect 1665 300 1695 326
rect 1761 300 1791 331
rect 1857 300 1887 326
rect 1953 300 1983 331
rect -1983 -331 -1953 -300
rect -1887 -326 -1857 -300
rect -1791 -331 -1761 -300
rect -1695 -326 -1665 -300
rect -1599 -331 -1569 -300
rect -1503 -326 -1473 -300
rect -1407 -331 -1377 -300
rect -1311 -326 -1281 -300
rect -1215 -331 -1185 -300
rect -1119 -326 -1089 -300
rect -1023 -331 -993 -300
rect -927 -326 -897 -300
rect -831 -331 -801 -300
rect -735 -326 -705 -300
rect -639 -331 -609 -300
rect -543 -326 -513 -300
rect -447 -331 -417 -300
rect -351 -326 -321 -300
rect -255 -331 -225 -300
rect -159 -326 -129 -300
rect -63 -331 -33 -300
rect 33 -326 63 -300
rect 129 -331 159 -300
rect 225 -326 255 -300
rect 321 -331 351 -300
rect 417 -326 447 -300
rect 513 -331 543 -300
rect 609 -326 639 -300
rect 705 -331 735 -300
rect 801 -326 831 -300
rect 897 -331 927 -300
rect 993 -326 1023 -300
rect 1089 -331 1119 -300
rect 1185 -326 1215 -300
rect 1281 -331 1311 -300
rect 1377 -326 1407 -300
rect 1473 -331 1503 -300
rect 1569 -326 1599 -300
rect 1665 -331 1695 -300
rect 1761 -326 1791 -300
rect 1857 -331 1887 -300
rect 1953 -326 1983 -300
rect -2001 -347 -1935 -331
rect -2001 -381 -1985 -347
rect -1951 -381 -1935 -347
rect -2001 -397 -1935 -381
rect -1809 -347 -1743 -331
rect -1809 -381 -1793 -347
rect -1759 -381 -1743 -347
rect -1809 -397 -1743 -381
rect -1617 -347 -1551 -331
rect -1617 -381 -1601 -347
rect -1567 -381 -1551 -347
rect -1617 -397 -1551 -381
rect -1425 -347 -1359 -331
rect -1425 -381 -1409 -347
rect -1375 -381 -1359 -347
rect -1425 -397 -1359 -381
rect -1233 -347 -1167 -331
rect -1233 -381 -1217 -347
rect -1183 -381 -1167 -347
rect -1233 -397 -1167 -381
rect -1041 -347 -975 -331
rect -1041 -381 -1025 -347
rect -991 -381 -975 -347
rect -1041 -397 -975 -381
rect -849 -347 -783 -331
rect -849 -381 -833 -347
rect -799 -381 -783 -347
rect -849 -397 -783 -381
rect -657 -347 -591 -331
rect -657 -381 -641 -347
rect -607 -381 -591 -347
rect -657 -397 -591 -381
rect -465 -347 -399 -331
rect -465 -381 -449 -347
rect -415 -381 -399 -347
rect -465 -397 -399 -381
rect -273 -347 -207 -331
rect -273 -381 -257 -347
rect -223 -381 -207 -347
rect -273 -397 -207 -381
rect -81 -347 -15 -331
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect -81 -397 -15 -381
rect 111 -347 177 -331
rect 111 -381 127 -347
rect 161 -381 177 -347
rect 111 -397 177 -381
rect 303 -347 369 -331
rect 303 -381 319 -347
rect 353 -381 369 -347
rect 303 -397 369 -381
rect 495 -347 561 -331
rect 495 -381 511 -347
rect 545 -381 561 -347
rect 495 -397 561 -381
rect 687 -347 753 -331
rect 687 -381 703 -347
rect 737 -381 753 -347
rect 687 -397 753 -381
rect 879 -347 945 -331
rect 879 -381 895 -347
rect 929 -381 945 -347
rect 879 -397 945 -381
rect 1071 -347 1137 -331
rect 1071 -381 1087 -347
rect 1121 -381 1137 -347
rect 1071 -397 1137 -381
rect 1263 -347 1329 -331
rect 1263 -381 1279 -347
rect 1313 -381 1329 -347
rect 1263 -397 1329 -381
rect 1455 -347 1521 -331
rect 1455 -381 1471 -347
rect 1505 -381 1521 -347
rect 1455 -397 1521 -381
rect 1647 -347 1713 -331
rect 1647 -381 1663 -347
rect 1697 -381 1713 -347
rect 1647 -397 1713 -381
rect 1839 -347 1905 -331
rect 1839 -381 1855 -347
rect 1889 -381 1905 -347
rect 1839 -397 1905 -381
<< polycont >>
rect -1889 347 -1855 381
rect -1697 347 -1663 381
rect -1505 347 -1471 381
rect -1313 347 -1279 381
rect -1121 347 -1087 381
rect -929 347 -895 381
rect -737 347 -703 381
rect -545 347 -511 381
rect -353 347 -319 381
rect -161 347 -127 381
rect 31 347 65 381
rect 223 347 257 381
rect 415 347 449 381
rect 607 347 641 381
rect 799 347 833 381
rect 991 347 1025 381
rect 1183 347 1217 381
rect 1375 347 1409 381
rect 1567 347 1601 381
rect 1759 347 1793 381
rect 1951 347 1985 381
rect -1985 -381 -1951 -347
rect -1793 -381 -1759 -347
rect -1601 -381 -1567 -347
rect -1409 -381 -1375 -347
rect -1217 -381 -1183 -347
rect -1025 -381 -991 -347
rect -833 -381 -799 -347
rect -641 -381 -607 -347
rect -449 -381 -415 -347
rect -257 -381 -223 -347
rect -65 -381 -31 -347
rect 127 -381 161 -347
rect 319 -381 353 -347
rect 511 -381 545 -347
rect 703 -381 737 -347
rect 895 -381 929 -347
rect 1087 -381 1121 -347
rect 1279 -381 1313 -347
rect 1471 -381 1505 -347
rect 1663 -381 1697 -347
rect 1855 -381 1889 -347
<< locali >>
rect -1905 347 -1889 381
rect -1855 347 -1839 381
rect -1713 347 -1697 381
rect -1663 347 -1647 381
rect -1521 347 -1505 381
rect -1471 347 -1455 381
rect -1329 347 -1313 381
rect -1279 347 -1263 381
rect -1137 347 -1121 381
rect -1087 347 -1071 381
rect -945 347 -929 381
rect -895 347 -879 381
rect -753 347 -737 381
rect -703 347 -687 381
rect -561 347 -545 381
rect -511 347 -495 381
rect -369 347 -353 381
rect -319 347 -303 381
rect -177 347 -161 381
rect -127 347 -111 381
rect 15 347 31 381
rect 65 347 81 381
rect 207 347 223 381
rect 257 347 273 381
rect 399 347 415 381
rect 449 347 465 381
rect 591 347 607 381
rect 641 347 657 381
rect 783 347 799 381
rect 833 347 849 381
rect 975 347 991 381
rect 1025 347 1041 381
rect 1167 347 1183 381
rect 1217 347 1233 381
rect 1359 347 1375 381
rect 1409 347 1425 381
rect 1551 347 1567 381
rect 1601 347 1617 381
rect 1743 347 1759 381
rect 1793 347 1809 381
rect 1935 347 1951 381
rect 1985 347 2001 381
rect -2033 269 -1999 304
rect -2033 197 -1999 221
rect -2033 125 -1999 153
rect -2033 53 -1999 85
rect -2033 -17 -1999 17
rect -2033 -85 -1999 -53
rect -2033 -153 -1999 -125
rect -2033 -221 -1999 -197
rect -2033 -304 -1999 -269
rect -1937 269 -1903 304
rect -1937 197 -1903 221
rect -1937 125 -1903 153
rect -1937 53 -1903 85
rect -1937 -17 -1903 17
rect -1937 -85 -1903 -53
rect -1937 -153 -1903 -125
rect -1937 -221 -1903 -197
rect -1937 -304 -1903 -269
rect -1841 269 -1807 304
rect -1841 197 -1807 221
rect -1841 125 -1807 153
rect -1841 53 -1807 85
rect -1841 -17 -1807 17
rect -1841 -85 -1807 -53
rect -1841 -153 -1807 -125
rect -1841 -221 -1807 -197
rect -1841 -304 -1807 -269
rect -1745 269 -1711 304
rect -1745 197 -1711 221
rect -1745 125 -1711 153
rect -1745 53 -1711 85
rect -1745 -17 -1711 17
rect -1745 -85 -1711 -53
rect -1745 -153 -1711 -125
rect -1745 -221 -1711 -197
rect -1745 -304 -1711 -269
rect -1649 269 -1615 304
rect -1649 197 -1615 221
rect -1649 125 -1615 153
rect -1649 53 -1615 85
rect -1649 -17 -1615 17
rect -1649 -85 -1615 -53
rect -1649 -153 -1615 -125
rect -1649 -221 -1615 -197
rect -1649 -304 -1615 -269
rect -1553 269 -1519 304
rect -1553 197 -1519 221
rect -1553 125 -1519 153
rect -1553 53 -1519 85
rect -1553 -17 -1519 17
rect -1553 -85 -1519 -53
rect -1553 -153 -1519 -125
rect -1553 -221 -1519 -197
rect -1553 -304 -1519 -269
rect -1457 269 -1423 304
rect -1457 197 -1423 221
rect -1457 125 -1423 153
rect -1457 53 -1423 85
rect -1457 -17 -1423 17
rect -1457 -85 -1423 -53
rect -1457 -153 -1423 -125
rect -1457 -221 -1423 -197
rect -1457 -304 -1423 -269
rect -1361 269 -1327 304
rect -1361 197 -1327 221
rect -1361 125 -1327 153
rect -1361 53 -1327 85
rect -1361 -17 -1327 17
rect -1361 -85 -1327 -53
rect -1361 -153 -1327 -125
rect -1361 -221 -1327 -197
rect -1361 -304 -1327 -269
rect -1265 269 -1231 304
rect -1265 197 -1231 221
rect -1265 125 -1231 153
rect -1265 53 -1231 85
rect -1265 -17 -1231 17
rect -1265 -85 -1231 -53
rect -1265 -153 -1231 -125
rect -1265 -221 -1231 -197
rect -1265 -304 -1231 -269
rect -1169 269 -1135 304
rect -1169 197 -1135 221
rect -1169 125 -1135 153
rect -1169 53 -1135 85
rect -1169 -17 -1135 17
rect -1169 -85 -1135 -53
rect -1169 -153 -1135 -125
rect -1169 -221 -1135 -197
rect -1169 -304 -1135 -269
rect -1073 269 -1039 304
rect -1073 197 -1039 221
rect -1073 125 -1039 153
rect -1073 53 -1039 85
rect -1073 -17 -1039 17
rect -1073 -85 -1039 -53
rect -1073 -153 -1039 -125
rect -1073 -221 -1039 -197
rect -1073 -304 -1039 -269
rect -977 269 -943 304
rect -977 197 -943 221
rect -977 125 -943 153
rect -977 53 -943 85
rect -977 -17 -943 17
rect -977 -85 -943 -53
rect -977 -153 -943 -125
rect -977 -221 -943 -197
rect -977 -304 -943 -269
rect -881 269 -847 304
rect -881 197 -847 221
rect -881 125 -847 153
rect -881 53 -847 85
rect -881 -17 -847 17
rect -881 -85 -847 -53
rect -881 -153 -847 -125
rect -881 -221 -847 -197
rect -881 -304 -847 -269
rect -785 269 -751 304
rect -785 197 -751 221
rect -785 125 -751 153
rect -785 53 -751 85
rect -785 -17 -751 17
rect -785 -85 -751 -53
rect -785 -153 -751 -125
rect -785 -221 -751 -197
rect -785 -304 -751 -269
rect -689 269 -655 304
rect -689 197 -655 221
rect -689 125 -655 153
rect -689 53 -655 85
rect -689 -17 -655 17
rect -689 -85 -655 -53
rect -689 -153 -655 -125
rect -689 -221 -655 -197
rect -689 -304 -655 -269
rect -593 269 -559 304
rect -593 197 -559 221
rect -593 125 -559 153
rect -593 53 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -53
rect -593 -153 -559 -125
rect -593 -221 -559 -197
rect -593 -304 -559 -269
rect -497 269 -463 304
rect -497 197 -463 221
rect -497 125 -463 153
rect -497 53 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -53
rect -497 -153 -463 -125
rect -497 -221 -463 -197
rect -497 -304 -463 -269
rect -401 269 -367 304
rect -401 197 -367 221
rect -401 125 -367 153
rect -401 53 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -53
rect -401 -153 -367 -125
rect -401 -221 -367 -197
rect -401 -304 -367 -269
rect -305 269 -271 304
rect -305 197 -271 221
rect -305 125 -271 153
rect -305 53 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -53
rect -305 -153 -271 -125
rect -305 -221 -271 -197
rect -305 -304 -271 -269
rect -209 269 -175 304
rect -209 197 -175 221
rect -209 125 -175 153
rect -209 53 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -53
rect -209 -153 -175 -125
rect -209 -221 -175 -197
rect -209 -304 -175 -269
rect -113 269 -79 304
rect -113 197 -79 221
rect -113 125 -79 153
rect -113 53 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -53
rect -113 -153 -79 -125
rect -113 -221 -79 -197
rect -113 -304 -79 -269
rect -17 269 17 304
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -304 17 -269
rect 79 269 113 304
rect 79 197 113 221
rect 79 125 113 153
rect 79 53 113 85
rect 79 -17 113 17
rect 79 -85 113 -53
rect 79 -153 113 -125
rect 79 -221 113 -197
rect 79 -304 113 -269
rect 175 269 209 304
rect 175 197 209 221
rect 175 125 209 153
rect 175 53 209 85
rect 175 -17 209 17
rect 175 -85 209 -53
rect 175 -153 209 -125
rect 175 -221 209 -197
rect 175 -304 209 -269
rect 271 269 305 304
rect 271 197 305 221
rect 271 125 305 153
rect 271 53 305 85
rect 271 -17 305 17
rect 271 -85 305 -53
rect 271 -153 305 -125
rect 271 -221 305 -197
rect 271 -304 305 -269
rect 367 269 401 304
rect 367 197 401 221
rect 367 125 401 153
rect 367 53 401 85
rect 367 -17 401 17
rect 367 -85 401 -53
rect 367 -153 401 -125
rect 367 -221 401 -197
rect 367 -304 401 -269
rect 463 269 497 304
rect 463 197 497 221
rect 463 125 497 153
rect 463 53 497 85
rect 463 -17 497 17
rect 463 -85 497 -53
rect 463 -153 497 -125
rect 463 -221 497 -197
rect 463 -304 497 -269
rect 559 269 593 304
rect 559 197 593 221
rect 559 125 593 153
rect 559 53 593 85
rect 559 -17 593 17
rect 559 -85 593 -53
rect 559 -153 593 -125
rect 559 -221 593 -197
rect 559 -304 593 -269
rect 655 269 689 304
rect 655 197 689 221
rect 655 125 689 153
rect 655 53 689 85
rect 655 -17 689 17
rect 655 -85 689 -53
rect 655 -153 689 -125
rect 655 -221 689 -197
rect 655 -304 689 -269
rect 751 269 785 304
rect 751 197 785 221
rect 751 125 785 153
rect 751 53 785 85
rect 751 -17 785 17
rect 751 -85 785 -53
rect 751 -153 785 -125
rect 751 -221 785 -197
rect 751 -304 785 -269
rect 847 269 881 304
rect 847 197 881 221
rect 847 125 881 153
rect 847 53 881 85
rect 847 -17 881 17
rect 847 -85 881 -53
rect 847 -153 881 -125
rect 847 -221 881 -197
rect 847 -304 881 -269
rect 943 269 977 304
rect 943 197 977 221
rect 943 125 977 153
rect 943 53 977 85
rect 943 -17 977 17
rect 943 -85 977 -53
rect 943 -153 977 -125
rect 943 -221 977 -197
rect 943 -304 977 -269
rect 1039 269 1073 304
rect 1039 197 1073 221
rect 1039 125 1073 153
rect 1039 53 1073 85
rect 1039 -17 1073 17
rect 1039 -85 1073 -53
rect 1039 -153 1073 -125
rect 1039 -221 1073 -197
rect 1039 -304 1073 -269
rect 1135 269 1169 304
rect 1135 197 1169 221
rect 1135 125 1169 153
rect 1135 53 1169 85
rect 1135 -17 1169 17
rect 1135 -85 1169 -53
rect 1135 -153 1169 -125
rect 1135 -221 1169 -197
rect 1135 -304 1169 -269
rect 1231 269 1265 304
rect 1231 197 1265 221
rect 1231 125 1265 153
rect 1231 53 1265 85
rect 1231 -17 1265 17
rect 1231 -85 1265 -53
rect 1231 -153 1265 -125
rect 1231 -221 1265 -197
rect 1231 -304 1265 -269
rect 1327 269 1361 304
rect 1327 197 1361 221
rect 1327 125 1361 153
rect 1327 53 1361 85
rect 1327 -17 1361 17
rect 1327 -85 1361 -53
rect 1327 -153 1361 -125
rect 1327 -221 1361 -197
rect 1327 -304 1361 -269
rect 1423 269 1457 304
rect 1423 197 1457 221
rect 1423 125 1457 153
rect 1423 53 1457 85
rect 1423 -17 1457 17
rect 1423 -85 1457 -53
rect 1423 -153 1457 -125
rect 1423 -221 1457 -197
rect 1423 -304 1457 -269
rect 1519 269 1553 304
rect 1519 197 1553 221
rect 1519 125 1553 153
rect 1519 53 1553 85
rect 1519 -17 1553 17
rect 1519 -85 1553 -53
rect 1519 -153 1553 -125
rect 1519 -221 1553 -197
rect 1519 -304 1553 -269
rect 1615 269 1649 304
rect 1615 197 1649 221
rect 1615 125 1649 153
rect 1615 53 1649 85
rect 1615 -17 1649 17
rect 1615 -85 1649 -53
rect 1615 -153 1649 -125
rect 1615 -221 1649 -197
rect 1615 -304 1649 -269
rect 1711 269 1745 304
rect 1711 197 1745 221
rect 1711 125 1745 153
rect 1711 53 1745 85
rect 1711 -17 1745 17
rect 1711 -85 1745 -53
rect 1711 -153 1745 -125
rect 1711 -221 1745 -197
rect 1711 -304 1745 -269
rect 1807 269 1841 304
rect 1807 197 1841 221
rect 1807 125 1841 153
rect 1807 53 1841 85
rect 1807 -17 1841 17
rect 1807 -85 1841 -53
rect 1807 -153 1841 -125
rect 1807 -221 1841 -197
rect 1807 -304 1841 -269
rect 1903 269 1937 304
rect 1903 197 1937 221
rect 1903 125 1937 153
rect 1903 53 1937 85
rect 1903 -17 1937 17
rect 1903 -85 1937 -53
rect 1903 -153 1937 -125
rect 1903 -221 1937 -197
rect 1903 -304 1937 -269
rect 1999 269 2033 304
rect 1999 197 2033 221
rect 1999 125 2033 153
rect 1999 53 2033 85
rect 1999 -17 2033 17
rect 1999 -85 2033 -53
rect 1999 -153 2033 -125
rect 1999 -221 2033 -197
rect 1999 -304 2033 -269
rect -2001 -381 -1985 -347
rect -1951 -381 -1935 -347
rect -1809 -381 -1793 -347
rect -1759 -381 -1743 -347
rect -1617 -381 -1601 -347
rect -1567 -381 -1551 -347
rect -1425 -381 -1409 -347
rect -1375 -381 -1359 -347
rect -1233 -381 -1217 -347
rect -1183 -381 -1167 -347
rect -1041 -381 -1025 -347
rect -991 -381 -975 -347
rect -849 -381 -833 -347
rect -799 -381 -783 -347
rect -657 -381 -641 -347
rect -607 -381 -591 -347
rect -465 -381 -449 -347
rect -415 -381 -399 -347
rect -273 -381 -257 -347
rect -223 -381 -207 -347
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect 111 -381 127 -347
rect 161 -381 177 -347
rect 303 -381 319 -347
rect 353 -381 369 -347
rect 495 -381 511 -347
rect 545 -381 561 -347
rect 687 -381 703 -347
rect 737 -381 753 -347
rect 879 -381 895 -347
rect 929 -381 945 -347
rect 1071 -381 1087 -347
rect 1121 -381 1137 -347
rect 1263 -381 1279 -347
rect 1313 -381 1329 -347
rect 1455 -381 1471 -347
rect 1505 -381 1521 -347
rect 1647 -381 1663 -347
rect 1697 -381 1713 -347
rect 1839 -381 1855 -347
rect 1889 -381 1905 -347
<< viali >>
rect -1889 347 -1855 381
rect -1697 347 -1663 381
rect -1505 347 -1471 381
rect -1313 347 -1279 381
rect -1121 347 -1087 381
rect -929 347 -895 381
rect -737 347 -703 381
rect -545 347 -511 381
rect -353 347 -319 381
rect -161 347 -127 381
rect 31 347 65 381
rect 223 347 257 381
rect 415 347 449 381
rect 607 347 641 381
rect 799 347 833 381
rect 991 347 1025 381
rect 1183 347 1217 381
rect 1375 347 1409 381
rect 1567 347 1601 381
rect 1759 347 1793 381
rect 1951 347 1985 381
rect -2033 255 -1999 269
rect -2033 235 -1999 255
rect -2033 187 -1999 197
rect -2033 163 -1999 187
rect -2033 119 -1999 125
rect -2033 91 -1999 119
rect -2033 51 -1999 53
rect -2033 19 -1999 51
rect -2033 -51 -1999 -19
rect -2033 -53 -1999 -51
rect -2033 -119 -1999 -91
rect -2033 -125 -1999 -119
rect -2033 -187 -1999 -163
rect -2033 -197 -1999 -187
rect -2033 -255 -1999 -235
rect -2033 -269 -1999 -255
rect -1937 255 -1903 269
rect -1937 235 -1903 255
rect -1937 187 -1903 197
rect -1937 163 -1903 187
rect -1937 119 -1903 125
rect -1937 91 -1903 119
rect -1937 51 -1903 53
rect -1937 19 -1903 51
rect -1937 -51 -1903 -19
rect -1937 -53 -1903 -51
rect -1937 -119 -1903 -91
rect -1937 -125 -1903 -119
rect -1937 -187 -1903 -163
rect -1937 -197 -1903 -187
rect -1937 -255 -1903 -235
rect -1937 -269 -1903 -255
rect -1841 255 -1807 269
rect -1841 235 -1807 255
rect -1841 187 -1807 197
rect -1841 163 -1807 187
rect -1841 119 -1807 125
rect -1841 91 -1807 119
rect -1841 51 -1807 53
rect -1841 19 -1807 51
rect -1841 -51 -1807 -19
rect -1841 -53 -1807 -51
rect -1841 -119 -1807 -91
rect -1841 -125 -1807 -119
rect -1841 -187 -1807 -163
rect -1841 -197 -1807 -187
rect -1841 -255 -1807 -235
rect -1841 -269 -1807 -255
rect -1745 255 -1711 269
rect -1745 235 -1711 255
rect -1745 187 -1711 197
rect -1745 163 -1711 187
rect -1745 119 -1711 125
rect -1745 91 -1711 119
rect -1745 51 -1711 53
rect -1745 19 -1711 51
rect -1745 -51 -1711 -19
rect -1745 -53 -1711 -51
rect -1745 -119 -1711 -91
rect -1745 -125 -1711 -119
rect -1745 -187 -1711 -163
rect -1745 -197 -1711 -187
rect -1745 -255 -1711 -235
rect -1745 -269 -1711 -255
rect -1649 255 -1615 269
rect -1649 235 -1615 255
rect -1649 187 -1615 197
rect -1649 163 -1615 187
rect -1649 119 -1615 125
rect -1649 91 -1615 119
rect -1649 51 -1615 53
rect -1649 19 -1615 51
rect -1649 -51 -1615 -19
rect -1649 -53 -1615 -51
rect -1649 -119 -1615 -91
rect -1649 -125 -1615 -119
rect -1649 -187 -1615 -163
rect -1649 -197 -1615 -187
rect -1649 -255 -1615 -235
rect -1649 -269 -1615 -255
rect -1553 255 -1519 269
rect -1553 235 -1519 255
rect -1553 187 -1519 197
rect -1553 163 -1519 187
rect -1553 119 -1519 125
rect -1553 91 -1519 119
rect -1553 51 -1519 53
rect -1553 19 -1519 51
rect -1553 -51 -1519 -19
rect -1553 -53 -1519 -51
rect -1553 -119 -1519 -91
rect -1553 -125 -1519 -119
rect -1553 -187 -1519 -163
rect -1553 -197 -1519 -187
rect -1553 -255 -1519 -235
rect -1553 -269 -1519 -255
rect -1457 255 -1423 269
rect -1457 235 -1423 255
rect -1457 187 -1423 197
rect -1457 163 -1423 187
rect -1457 119 -1423 125
rect -1457 91 -1423 119
rect -1457 51 -1423 53
rect -1457 19 -1423 51
rect -1457 -51 -1423 -19
rect -1457 -53 -1423 -51
rect -1457 -119 -1423 -91
rect -1457 -125 -1423 -119
rect -1457 -187 -1423 -163
rect -1457 -197 -1423 -187
rect -1457 -255 -1423 -235
rect -1457 -269 -1423 -255
rect -1361 255 -1327 269
rect -1361 235 -1327 255
rect -1361 187 -1327 197
rect -1361 163 -1327 187
rect -1361 119 -1327 125
rect -1361 91 -1327 119
rect -1361 51 -1327 53
rect -1361 19 -1327 51
rect -1361 -51 -1327 -19
rect -1361 -53 -1327 -51
rect -1361 -119 -1327 -91
rect -1361 -125 -1327 -119
rect -1361 -187 -1327 -163
rect -1361 -197 -1327 -187
rect -1361 -255 -1327 -235
rect -1361 -269 -1327 -255
rect -1265 255 -1231 269
rect -1265 235 -1231 255
rect -1265 187 -1231 197
rect -1265 163 -1231 187
rect -1265 119 -1231 125
rect -1265 91 -1231 119
rect -1265 51 -1231 53
rect -1265 19 -1231 51
rect -1265 -51 -1231 -19
rect -1265 -53 -1231 -51
rect -1265 -119 -1231 -91
rect -1265 -125 -1231 -119
rect -1265 -187 -1231 -163
rect -1265 -197 -1231 -187
rect -1265 -255 -1231 -235
rect -1265 -269 -1231 -255
rect -1169 255 -1135 269
rect -1169 235 -1135 255
rect -1169 187 -1135 197
rect -1169 163 -1135 187
rect -1169 119 -1135 125
rect -1169 91 -1135 119
rect -1169 51 -1135 53
rect -1169 19 -1135 51
rect -1169 -51 -1135 -19
rect -1169 -53 -1135 -51
rect -1169 -119 -1135 -91
rect -1169 -125 -1135 -119
rect -1169 -187 -1135 -163
rect -1169 -197 -1135 -187
rect -1169 -255 -1135 -235
rect -1169 -269 -1135 -255
rect -1073 255 -1039 269
rect -1073 235 -1039 255
rect -1073 187 -1039 197
rect -1073 163 -1039 187
rect -1073 119 -1039 125
rect -1073 91 -1039 119
rect -1073 51 -1039 53
rect -1073 19 -1039 51
rect -1073 -51 -1039 -19
rect -1073 -53 -1039 -51
rect -1073 -119 -1039 -91
rect -1073 -125 -1039 -119
rect -1073 -187 -1039 -163
rect -1073 -197 -1039 -187
rect -1073 -255 -1039 -235
rect -1073 -269 -1039 -255
rect -977 255 -943 269
rect -977 235 -943 255
rect -977 187 -943 197
rect -977 163 -943 187
rect -977 119 -943 125
rect -977 91 -943 119
rect -977 51 -943 53
rect -977 19 -943 51
rect -977 -51 -943 -19
rect -977 -53 -943 -51
rect -977 -119 -943 -91
rect -977 -125 -943 -119
rect -977 -187 -943 -163
rect -977 -197 -943 -187
rect -977 -255 -943 -235
rect -977 -269 -943 -255
rect -881 255 -847 269
rect -881 235 -847 255
rect -881 187 -847 197
rect -881 163 -847 187
rect -881 119 -847 125
rect -881 91 -847 119
rect -881 51 -847 53
rect -881 19 -847 51
rect -881 -51 -847 -19
rect -881 -53 -847 -51
rect -881 -119 -847 -91
rect -881 -125 -847 -119
rect -881 -187 -847 -163
rect -881 -197 -847 -187
rect -881 -255 -847 -235
rect -881 -269 -847 -255
rect -785 255 -751 269
rect -785 235 -751 255
rect -785 187 -751 197
rect -785 163 -751 187
rect -785 119 -751 125
rect -785 91 -751 119
rect -785 51 -751 53
rect -785 19 -751 51
rect -785 -51 -751 -19
rect -785 -53 -751 -51
rect -785 -119 -751 -91
rect -785 -125 -751 -119
rect -785 -187 -751 -163
rect -785 -197 -751 -187
rect -785 -255 -751 -235
rect -785 -269 -751 -255
rect -689 255 -655 269
rect -689 235 -655 255
rect -689 187 -655 197
rect -689 163 -655 187
rect -689 119 -655 125
rect -689 91 -655 119
rect -689 51 -655 53
rect -689 19 -655 51
rect -689 -51 -655 -19
rect -689 -53 -655 -51
rect -689 -119 -655 -91
rect -689 -125 -655 -119
rect -689 -187 -655 -163
rect -689 -197 -655 -187
rect -689 -255 -655 -235
rect -689 -269 -655 -255
rect -593 255 -559 269
rect -593 235 -559 255
rect -593 187 -559 197
rect -593 163 -559 187
rect -593 119 -559 125
rect -593 91 -559 119
rect -593 51 -559 53
rect -593 19 -559 51
rect -593 -51 -559 -19
rect -593 -53 -559 -51
rect -593 -119 -559 -91
rect -593 -125 -559 -119
rect -593 -187 -559 -163
rect -593 -197 -559 -187
rect -593 -255 -559 -235
rect -593 -269 -559 -255
rect -497 255 -463 269
rect -497 235 -463 255
rect -497 187 -463 197
rect -497 163 -463 187
rect -497 119 -463 125
rect -497 91 -463 119
rect -497 51 -463 53
rect -497 19 -463 51
rect -497 -51 -463 -19
rect -497 -53 -463 -51
rect -497 -119 -463 -91
rect -497 -125 -463 -119
rect -497 -187 -463 -163
rect -497 -197 -463 -187
rect -497 -255 -463 -235
rect -497 -269 -463 -255
rect -401 255 -367 269
rect -401 235 -367 255
rect -401 187 -367 197
rect -401 163 -367 187
rect -401 119 -367 125
rect -401 91 -367 119
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -401 -119 -367 -91
rect -401 -125 -367 -119
rect -401 -187 -367 -163
rect -401 -197 -367 -187
rect -401 -255 -367 -235
rect -401 -269 -367 -255
rect -305 255 -271 269
rect -305 235 -271 255
rect -305 187 -271 197
rect -305 163 -271 187
rect -305 119 -271 125
rect -305 91 -271 119
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -305 -119 -271 -91
rect -305 -125 -271 -119
rect -305 -187 -271 -163
rect -305 -197 -271 -187
rect -305 -255 -271 -235
rect -305 -269 -271 -255
rect -209 255 -175 269
rect -209 235 -175 255
rect -209 187 -175 197
rect -209 163 -175 187
rect -209 119 -175 125
rect -209 91 -175 119
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -209 -119 -175 -91
rect -209 -125 -175 -119
rect -209 -187 -175 -163
rect -209 -197 -175 -187
rect -209 -255 -175 -235
rect -209 -269 -175 -255
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 175 255 209 269
rect 175 235 209 255
rect 175 187 209 197
rect 175 163 209 187
rect 175 119 209 125
rect 175 91 209 119
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 175 -119 209 -91
rect 175 -125 209 -119
rect 175 -187 209 -163
rect 175 -197 209 -187
rect 175 -255 209 -235
rect 175 -269 209 -255
rect 271 255 305 269
rect 271 235 305 255
rect 271 187 305 197
rect 271 163 305 187
rect 271 119 305 125
rect 271 91 305 119
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect 271 -119 305 -91
rect 271 -125 305 -119
rect 271 -187 305 -163
rect 271 -197 305 -187
rect 271 -255 305 -235
rect 271 -269 305 -255
rect 367 255 401 269
rect 367 235 401 255
rect 367 187 401 197
rect 367 163 401 187
rect 367 119 401 125
rect 367 91 401 119
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 367 -119 401 -91
rect 367 -125 401 -119
rect 367 -187 401 -163
rect 367 -197 401 -187
rect 367 -255 401 -235
rect 367 -269 401 -255
rect 463 255 497 269
rect 463 235 497 255
rect 463 187 497 197
rect 463 163 497 187
rect 463 119 497 125
rect 463 91 497 119
rect 463 51 497 53
rect 463 19 497 51
rect 463 -51 497 -19
rect 463 -53 497 -51
rect 463 -119 497 -91
rect 463 -125 497 -119
rect 463 -187 497 -163
rect 463 -197 497 -187
rect 463 -255 497 -235
rect 463 -269 497 -255
rect 559 255 593 269
rect 559 235 593 255
rect 559 187 593 197
rect 559 163 593 187
rect 559 119 593 125
rect 559 91 593 119
rect 559 51 593 53
rect 559 19 593 51
rect 559 -51 593 -19
rect 559 -53 593 -51
rect 559 -119 593 -91
rect 559 -125 593 -119
rect 559 -187 593 -163
rect 559 -197 593 -187
rect 559 -255 593 -235
rect 559 -269 593 -255
rect 655 255 689 269
rect 655 235 689 255
rect 655 187 689 197
rect 655 163 689 187
rect 655 119 689 125
rect 655 91 689 119
rect 655 51 689 53
rect 655 19 689 51
rect 655 -51 689 -19
rect 655 -53 689 -51
rect 655 -119 689 -91
rect 655 -125 689 -119
rect 655 -187 689 -163
rect 655 -197 689 -187
rect 655 -255 689 -235
rect 655 -269 689 -255
rect 751 255 785 269
rect 751 235 785 255
rect 751 187 785 197
rect 751 163 785 187
rect 751 119 785 125
rect 751 91 785 119
rect 751 51 785 53
rect 751 19 785 51
rect 751 -51 785 -19
rect 751 -53 785 -51
rect 751 -119 785 -91
rect 751 -125 785 -119
rect 751 -187 785 -163
rect 751 -197 785 -187
rect 751 -255 785 -235
rect 751 -269 785 -255
rect 847 255 881 269
rect 847 235 881 255
rect 847 187 881 197
rect 847 163 881 187
rect 847 119 881 125
rect 847 91 881 119
rect 847 51 881 53
rect 847 19 881 51
rect 847 -51 881 -19
rect 847 -53 881 -51
rect 847 -119 881 -91
rect 847 -125 881 -119
rect 847 -187 881 -163
rect 847 -197 881 -187
rect 847 -255 881 -235
rect 847 -269 881 -255
rect 943 255 977 269
rect 943 235 977 255
rect 943 187 977 197
rect 943 163 977 187
rect 943 119 977 125
rect 943 91 977 119
rect 943 51 977 53
rect 943 19 977 51
rect 943 -51 977 -19
rect 943 -53 977 -51
rect 943 -119 977 -91
rect 943 -125 977 -119
rect 943 -187 977 -163
rect 943 -197 977 -187
rect 943 -255 977 -235
rect 943 -269 977 -255
rect 1039 255 1073 269
rect 1039 235 1073 255
rect 1039 187 1073 197
rect 1039 163 1073 187
rect 1039 119 1073 125
rect 1039 91 1073 119
rect 1039 51 1073 53
rect 1039 19 1073 51
rect 1039 -51 1073 -19
rect 1039 -53 1073 -51
rect 1039 -119 1073 -91
rect 1039 -125 1073 -119
rect 1039 -187 1073 -163
rect 1039 -197 1073 -187
rect 1039 -255 1073 -235
rect 1039 -269 1073 -255
rect 1135 255 1169 269
rect 1135 235 1169 255
rect 1135 187 1169 197
rect 1135 163 1169 187
rect 1135 119 1169 125
rect 1135 91 1169 119
rect 1135 51 1169 53
rect 1135 19 1169 51
rect 1135 -51 1169 -19
rect 1135 -53 1169 -51
rect 1135 -119 1169 -91
rect 1135 -125 1169 -119
rect 1135 -187 1169 -163
rect 1135 -197 1169 -187
rect 1135 -255 1169 -235
rect 1135 -269 1169 -255
rect 1231 255 1265 269
rect 1231 235 1265 255
rect 1231 187 1265 197
rect 1231 163 1265 187
rect 1231 119 1265 125
rect 1231 91 1265 119
rect 1231 51 1265 53
rect 1231 19 1265 51
rect 1231 -51 1265 -19
rect 1231 -53 1265 -51
rect 1231 -119 1265 -91
rect 1231 -125 1265 -119
rect 1231 -187 1265 -163
rect 1231 -197 1265 -187
rect 1231 -255 1265 -235
rect 1231 -269 1265 -255
rect 1327 255 1361 269
rect 1327 235 1361 255
rect 1327 187 1361 197
rect 1327 163 1361 187
rect 1327 119 1361 125
rect 1327 91 1361 119
rect 1327 51 1361 53
rect 1327 19 1361 51
rect 1327 -51 1361 -19
rect 1327 -53 1361 -51
rect 1327 -119 1361 -91
rect 1327 -125 1361 -119
rect 1327 -187 1361 -163
rect 1327 -197 1361 -187
rect 1327 -255 1361 -235
rect 1327 -269 1361 -255
rect 1423 255 1457 269
rect 1423 235 1457 255
rect 1423 187 1457 197
rect 1423 163 1457 187
rect 1423 119 1457 125
rect 1423 91 1457 119
rect 1423 51 1457 53
rect 1423 19 1457 51
rect 1423 -51 1457 -19
rect 1423 -53 1457 -51
rect 1423 -119 1457 -91
rect 1423 -125 1457 -119
rect 1423 -187 1457 -163
rect 1423 -197 1457 -187
rect 1423 -255 1457 -235
rect 1423 -269 1457 -255
rect 1519 255 1553 269
rect 1519 235 1553 255
rect 1519 187 1553 197
rect 1519 163 1553 187
rect 1519 119 1553 125
rect 1519 91 1553 119
rect 1519 51 1553 53
rect 1519 19 1553 51
rect 1519 -51 1553 -19
rect 1519 -53 1553 -51
rect 1519 -119 1553 -91
rect 1519 -125 1553 -119
rect 1519 -187 1553 -163
rect 1519 -197 1553 -187
rect 1519 -255 1553 -235
rect 1519 -269 1553 -255
rect 1615 255 1649 269
rect 1615 235 1649 255
rect 1615 187 1649 197
rect 1615 163 1649 187
rect 1615 119 1649 125
rect 1615 91 1649 119
rect 1615 51 1649 53
rect 1615 19 1649 51
rect 1615 -51 1649 -19
rect 1615 -53 1649 -51
rect 1615 -119 1649 -91
rect 1615 -125 1649 -119
rect 1615 -187 1649 -163
rect 1615 -197 1649 -187
rect 1615 -255 1649 -235
rect 1615 -269 1649 -255
rect 1711 255 1745 269
rect 1711 235 1745 255
rect 1711 187 1745 197
rect 1711 163 1745 187
rect 1711 119 1745 125
rect 1711 91 1745 119
rect 1711 51 1745 53
rect 1711 19 1745 51
rect 1711 -51 1745 -19
rect 1711 -53 1745 -51
rect 1711 -119 1745 -91
rect 1711 -125 1745 -119
rect 1711 -187 1745 -163
rect 1711 -197 1745 -187
rect 1711 -255 1745 -235
rect 1711 -269 1745 -255
rect 1807 255 1841 269
rect 1807 235 1841 255
rect 1807 187 1841 197
rect 1807 163 1841 187
rect 1807 119 1841 125
rect 1807 91 1841 119
rect 1807 51 1841 53
rect 1807 19 1841 51
rect 1807 -51 1841 -19
rect 1807 -53 1841 -51
rect 1807 -119 1841 -91
rect 1807 -125 1841 -119
rect 1807 -187 1841 -163
rect 1807 -197 1841 -187
rect 1807 -255 1841 -235
rect 1807 -269 1841 -255
rect 1903 255 1937 269
rect 1903 235 1937 255
rect 1903 187 1937 197
rect 1903 163 1937 187
rect 1903 119 1937 125
rect 1903 91 1937 119
rect 1903 51 1937 53
rect 1903 19 1937 51
rect 1903 -51 1937 -19
rect 1903 -53 1937 -51
rect 1903 -119 1937 -91
rect 1903 -125 1937 -119
rect 1903 -187 1937 -163
rect 1903 -197 1937 -187
rect 1903 -255 1937 -235
rect 1903 -269 1937 -255
rect 1999 255 2033 269
rect 1999 235 2033 255
rect 1999 187 2033 197
rect 1999 163 2033 187
rect 1999 119 2033 125
rect 1999 91 2033 119
rect 1999 51 2033 53
rect 1999 19 2033 51
rect 1999 -51 2033 -19
rect 1999 -53 2033 -51
rect 1999 -119 2033 -91
rect 1999 -125 2033 -119
rect 1999 -187 2033 -163
rect 1999 -197 2033 -187
rect 1999 -255 2033 -235
rect 1999 -269 2033 -255
rect -1985 -381 -1951 -347
rect -1793 -381 -1759 -347
rect -1601 -381 -1567 -347
rect -1409 -381 -1375 -347
rect -1217 -381 -1183 -347
rect -1025 -381 -991 -347
rect -833 -381 -799 -347
rect -641 -381 -607 -347
rect -449 -381 -415 -347
rect -257 -381 -223 -347
rect -65 -381 -31 -347
rect 127 -381 161 -347
rect 319 -381 353 -347
rect 511 -381 545 -347
rect 703 -381 737 -347
rect 895 -381 929 -347
rect 1087 -381 1121 -347
rect 1279 -381 1313 -347
rect 1471 -381 1505 -347
rect 1663 -381 1697 -347
rect 1855 -381 1889 -347
<< metal1 >>
rect -1901 381 -1843 387
rect -1901 347 -1889 381
rect -1855 347 -1843 381
rect -1901 341 -1843 347
rect -1709 381 -1651 387
rect -1709 347 -1697 381
rect -1663 347 -1651 381
rect -1709 341 -1651 347
rect -1517 381 -1459 387
rect -1517 347 -1505 381
rect -1471 347 -1459 381
rect -1517 341 -1459 347
rect -1325 381 -1267 387
rect -1325 347 -1313 381
rect -1279 347 -1267 381
rect -1325 341 -1267 347
rect -1133 381 -1075 387
rect -1133 347 -1121 381
rect -1087 347 -1075 381
rect -1133 341 -1075 347
rect -941 381 -883 387
rect -941 347 -929 381
rect -895 347 -883 381
rect -941 341 -883 347
rect -749 381 -691 387
rect -749 347 -737 381
rect -703 347 -691 381
rect -749 341 -691 347
rect -557 381 -499 387
rect -557 347 -545 381
rect -511 347 -499 381
rect -557 341 -499 347
rect -365 381 -307 387
rect -365 347 -353 381
rect -319 347 -307 381
rect -365 341 -307 347
rect -173 381 -115 387
rect -173 347 -161 381
rect -127 347 -115 381
rect -173 341 -115 347
rect 19 381 77 387
rect 19 347 31 381
rect 65 347 77 381
rect 19 341 77 347
rect 211 381 269 387
rect 211 347 223 381
rect 257 347 269 381
rect 211 341 269 347
rect 403 381 461 387
rect 403 347 415 381
rect 449 347 461 381
rect 403 341 461 347
rect 595 381 653 387
rect 595 347 607 381
rect 641 347 653 381
rect 595 341 653 347
rect 787 381 845 387
rect 787 347 799 381
rect 833 347 845 381
rect 787 341 845 347
rect 979 381 1037 387
rect 979 347 991 381
rect 1025 347 1037 381
rect 979 341 1037 347
rect 1171 381 1229 387
rect 1171 347 1183 381
rect 1217 347 1229 381
rect 1171 341 1229 347
rect 1363 381 1421 387
rect 1363 347 1375 381
rect 1409 347 1421 381
rect 1363 341 1421 347
rect 1555 381 1613 387
rect 1555 347 1567 381
rect 1601 347 1613 381
rect 1555 341 1613 347
rect 1747 381 1805 387
rect 1747 347 1759 381
rect 1793 347 1805 381
rect 1747 341 1805 347
rect 1939 381 1997 387
rect 1939 347 1951 381
rect 1985 347 1997 381
rect 1939 341 1997 347
rect -2039 269 -1993 300
rect -2039 235 -2033 269
rect -1999 235 -1993 269
rect -2039 197 -1993 235
rect -2039 163 -2033 197
rect -1999 163 -1993 197
rect -2039 125 -1993 163
rect -2039 91 -2033 125
rect -1999 91 -1993 125
rect -2039 53 -1993 91
rect -2039 19 -2033 53
rect -1999 19 -1993 53
rect -2039 -19 -1993 19
rect -2039 -53 -2033 -19
rect -1999 -53 -1993 -19
rect -2039 -91 -1993 -53
rect -2039 -125 -2033 -91
rect -1999 -125 -1993 -91
rect -2039 -163 -1993 -125
rect -2039 -197 -2033 -163
rect -1999 -197 -1993 -163
rect -2039 -235 -1993 -197
rect -2039 -269 -2033 -235
rect -1999 -269 -1993 -235
rect -2039 -300 -1993 -269
rect -1943 269 -1897 300
rect -1943 235 -1937 269
rect -1903 235 -1897 269
rect -1943 197 -1897 235
rect -1943 163 -1937 197
rect -1903 163 -1897 197
rect -1943 125 -1897 163
rect -1943 91 -1937 125
rect -1903 91 -1897 125
rect -1943 53 -1897 91
rect -1943 19 -1937 53
rect -1903 19 -1897 53
rect -1943 -19 -1897 19
rect -1943 -53 -1937 -19
rect -1903 -53 -1897 -19
rect -1943 -91 -1897 -53
rect -1943 -125 -1937 -91
rect -1903 -125 -1897 -91
rect -1943 -163 -1897 -125
rect -1943 -197 -1937 -163
rect -1903 -197 -1897 -163
rect -1943 -235 -1897 -197
rect -1943 -269 -1937 -235
rect -1903 -269 -1897 -235
rect -1943 -300 -1897 -269
rect -1847 269 -1801 300
rect -1847 235 -1841 269
rect -1807 235 -1801 269
rect -1847 197 -1801 235
rect -1847 163 -1841 197
rect -1807 163 -1801 197
rect -1847 125 -1801 163
rect -1847 91 -1841 125
rect -1807 91 -1801 125
rect -1847 53 -1801 91
rect -1847 19 -1841 53
rect -1807 19 -1801 53
rect -1847 -19 -1801 19
rect -1847 -53 -1841 -19
rect -1807 -53 -1801 -19
rect -1847 -91 -1801 -53
rect -1847 -125 -1841 -91
rect -1807 -125 -1801 -91
rect -1847 -163 -1801 -125
rect -1847 -197 -1841 -163
rect -1807 -197 -1801 -163
rect -1847 -235 -1801 -197
rect -1847 -269 -1841 -235
rect -1807 -269 -1801 -235
rect -1847 -300 -1801 -269
rect -1751 269 -1705 300
rect -1751 235 -1745 269
rect -1711 235 -1705 269
rect -1751 197 -1705 235
rect -1751 163 -1745 197
rect -1711 163 -1705 197
rect -1751 125 -1705 163
rect -1751 91 -1745 125
rect -1711 91 -1705 125
rect -1751 53 -1705 91
rect -1751 19 -1745 53
rect -1711 19 -1705 53
rect -1751 -19 -1705 19
rect -1751 -53 -1745 -19
rect -1711 -53 -1705 -19
rect -1751 -91 -1705 -53
rect -1751 -125 -1745 -91
rect -1711 -125 -1705 -91
rect -1751 -163 -1705 -125
rect -1751 -197 -1745 -163
rect -1711 -197 -1705 -163
rect -1751 -235 -1705 -197
rect -1751 -269 -1745 -235
rect -1711 -269 -1705 -235
rect -1751 -300 -1705 -269
rect -1655 269 -1609 300
rect -1655 235 -1649 269
rect -1615 235 -1609 269
rect -1655 197 -1609 235
rect -1655 163 -1649 197
rect -1615 163 -1609 197
rect -1655 125 -1609 163
rect -1655 91 -1649 125
rect -1615 91 -1609 125
rect -1655 53 -1609 91
rect -1655 19 -1649 53
rect -1615 19 -1609 53
rect -1655 -19 -1609 19
rect -1655 -53 -1649 -19
rect -1615 -53 -1609 -19
rect -1655 -91 -1609 -53
rect -1655 -125 -1649 -91
rect -1615 -125 -1609 -91
rect -1655 -163 -1609 -125
rect -1655 -197 -1649 -163
rect -1615 -197 -1609 -163
rect -1655 -235 -1609 -197
rect -1655 -269 -1649 -235
rect -1615 -269 -1609 -235
rect -1655 -300 -1609 -269
rect -1559 269 -1513 300
rect -1559 235 -1553 269
rect -1519 235 -1513 269
rect -1559 197 -1513 235
rect -1559 163 -1553 197
rect -1519 163 -1513 197
rect -1559 125 -1513 163
rect -1559 91 -1553 125
rect -1519 91 -1513 125
rect -1559 53 -1513 91
rect -1559 19 -1553 53
rect -1519 19 -1513 53
rect -1559 -19 -1513 19
rect -1559 -53 -1553 -19
rect -1519 -53 -1513 -19
rect -1559 -91 -1513 -53
rect -1559 -125 -1553 -91
rect -1519 -125 -1513 -91
rect -1559 -163 -1513 -125
rect -1559 -197 -1553 -163
rect -1519 -197 -1513 -163
rect -1559 -235 -1513 -197
rect -1559 -269 -1553 -235
rect -1519 -269 -1513 -235
rect -1559 -300 -1513 -269
rect -1463 269 -1417 300
rect -1463 235 -1457 269
rect -1423 235 -1417 269
rect -1463 197 -1417 235
rect -1463 163 -1457 197
rect -1423 163 -1417 197
rect -1463 125 -1417 163
rect -1463 91 -1457 125
rect -1423 91 -1417 125
rect -1463 53 -1417 91
rect -1463 19 -1457 53
rect -1423 19 -1417 53
rect -1463 -19 -1417 19
rect -1463 -53 -1457 -19
rect -1423 -53 -1417 -19
rect -1463 -91 -1417 -53
rect -1463 -125 -1457 -91
rect -1423 -125 -1417 -91
rect -1463 -163 -1417 -125
rect -1463 -197 -1457 -163
rect -1423 -197 -1417 -163
rect -1463 -235 -1417 -197
rect -1463 -269 -1457 -235
rect -1423 -269 -1417 -235
rect -1463 -300 -1417 -269
rect -1367 269 -1321 300
rect -1367 235 -1361 269
rect -1327 235 -1321 269
rect -1367 197 -1321 235
rect -1367 163 -1361 197
rect -1327 163 -1321 197
rect -1367 125 -1321 163
rect -1367 91 -1361 125
rect -1327 91 -1321 125
rect -1367 53 -1321 91
rect -1367 19 -1361 53
rect -1327 19 -1321 53
rect -1367 -19 -1321 19
rect -1367 -53 -1361 -19
rect -1327 -53 -1321 -19
rect -1367 -91 -1321 -53
rect -1367 -125 -1361 -91
rect -1327 -125 -1321 -91
rect -1367 -163 -1321 -125
rect -1367 -197 -1361 -163
rect -1327 -197 -1321 -163
rect -1367 -235 -1321 -197
rect -1367 -269 -1361 -235
rect -1327 -269 -1321 -235
rect -1367 -300 -1321 -269
rect -1271 269 -1225 300
rect -1271 235 -1265 269
rect -1231 235 -1225 269
rect -1271 197 -1225 235
rect -1271 163 -1265 197
rect -1231 163 -1225 197
rect -1271 125 -1225 163
rect -1271 91 -1265 125
rect -1231 91 -1225 125
rect -1271 53 -1225 91
rect -1271 19 -1265 53
rect -1231 19 -1225 53
rect -1271 -19 -1225 19
rect -1271 -53 -1265 -19
rect -1231 -53 -1225 -19
rect -1271 -91 -1225 -53
rect -1271 -125 -1265 -91
rect -1231 -125 -1225 -91
rect -1271 -163 -1225 -125
rect -1271 -197 -1265 -163
rect -1231 -197 -1225 -163
rect -1271 -235 -1225 -197
rect -1271 -269 -1265 -235
rect -1231 -269 -1225 -235
rect -1271 -300 -1225 -269
rect -1175 269 -1129 300
rect -1175 235 -1169 269
rect -1135 235 -1129 269
rect -1175 197 -1129 235
rect -1175 163 -1169 197
rect -1135 163 -1129 197
rect -1175 125 -1129 163
rect -1175 91 -1169 125
rect -1135 91 -1129 125
rect -1175 53 -1129 91
rect -1175 19 -1169 53
rect -1135 19 -1129 53
rect -1175 -19 -1129 19
rect -1175 -53 -1169 -19
rect -1135 -53 -1129 -19
rect -1175 -91 -1129 -53
rect -1175 -125 -1169 -91
rect -1135 -125 -1129 -91
rect -1175 -163 -1129 -125
rect -1175 -197 -1169 -163
rect -1135 -197 -1129 -163
rect -1175 -235 -1129 -197
rect -1175 -269 -1169 -235
rect -1135 -269 -1129 -235
rect -1175 -300 -1129 -269
rect -1079 269 -1033 300
rect -1079 235 -1073 269
rect -1039 235 -1033 269
rect -1079 197 -1033 235
rect -1079 163 -1073 197
rect -1039 163 -1033 197
rect -1079 125 -1033 163
rect -1079 91 -1073 125
rect -1039 91 -1033 125
rect -1079 53 -1033 91
rect -1079 19 -1073 53
rect -1039 19 -1033 53
rect -1079 -19 -1033 19
rect -1079 -53 -1073 -19
rect -1039 -53 -1033 -19
rect -1079 -91 -1033 -53
rect -1079 -125 -1073 -91
rect -1039 -125 -1033 -91
rect -1079 -163 -1033 -125
rect -1079 -197 -1073 -163
rect -1039 -197 -1033 -163
rect -1079 -235 -1033 -197
rect -1079 -269 -1073 -235
rect -1039 -269 -1033 -235
rect -1079 -300 -1033 -269
rect -983 269 -937 300
rect -983 235 -977 269
rect -943 235 -937 269
rect -983 197 -937 235
rect -983 163 -977 197
rect -943 163 -937 197
rect -983 125 -937 163
rect -983 91 -977 125
rect -943 91 -937 125
rect -983 53 -937 91
rect -983 19 -977 53
rect -943 19 -937 53
rect -983 -19 -937 19
rect -983 -53 -977 -19
rect -943 -53 -937 -19
rect -983 -91 -937 -53
rect -983 -125 -977 -91
rect -943 -125 -937 -91
rect -983 -163 -937 -125
rect -983 -197 -977 -163
rect -943 -197 -937 -163
rect -983 -235 -937 -197
rect -983 -269 -977 -235
rect -943 -269 -937 -235
rect -983 -300 -937 -269
rect -887 269 -841 300
rect -887 235 -881 269
rect -847 235 -841 269
rect -887 197 -841 235
rect -887 163 -881 197
rect -847 163 -841 197
rect -887 125 -841 163
rect -887 91 -881 125
rect -847 91 -841 125
rect -887 53 -841 91
rect -887 19 -881 53
rect -847 19 -841 53
rect -887 -19 -841 19
rect -887 -53 -881 -19
rect -847 -53 -841 -19
rect -887 -91 -841 -53
rect -887 -125 -881 -91
rect -847 -125 -841 -91
rect -887 -163 -841 -125
rect -887 -197 -881 -163
rect -847 -197 -841 -163
rect -887 -235 -841 -197
rect -887 -269 -881 -235
rect -847 -269 -841 -235
rect -887 -300 -841 -269
rect -791 269 -745 300
rect -791 235 -785 269
rect -751 235 -745 269
rect -791 197 -745 235
rect -791 163 -785 197
rect -751 163 -745 197
rect -791 125 -745 163
rect -791 91 -785 125
rect -751 91 -745 125
rect -791 53 -745 91
rect -791 19 -785 53
rect -751 19 -745 53
rect -791 -19 -745 19
rect -791 -53 -785 -19
rect -751 -53 -745 -19
rect -791 -91 -745 -53
rect -791 -125 -785 -91
rect -751 -125 -745 -91
rect -791 -163 -745 -125
rect -791 -197 -785 -163
rect -751 -197 -745 -163
rect -791 -235 -745 -197
rect -791 -269 -785 -235
rect -751 -269 -745 -235
rect -791 -300 -745 -269
rect -695 269 -649 300
rect -695 235 -689 269
rect -655 235 -649 269
rect -695 197 -649 235
rect -695 163 -689 197
rect -655 163 -649 197
rect -695 125 -649 163
rect -695 91 -689 125
rect -655 91 -649 125
rect -695 53 -649 91
rect -695 19 -689 53
rect -655 19 -649 53
rect -695 -19 -649 19
rect -695 -53 -689 -19
rect -655 -53 -649 -19
rect -695 -91 -649 -53
rect -695 -125 -689 -91
rect -655 -125 -649 -91
rect -695 -163 -649 -125
rect -695 -197 -689 -163
rect -655 -197 -649 -163
rect -695 -235 -649 -197
rect -695 -269 -689 -235
rect -655 -269 -649 -235
rect -695 -300 -649 -269
rect -599 269 -553 300
rect -599 235 -593 269
rect -559 235 -553 269
rect -599 197 -553 235
rect -599 163 -593 197
rect -559 163 -553 197
rect -599 125 -553 163
rect -599 91 -593 125
rect -559 91 -553 125
rect -599 53 -553 91
rect -599 19 -593 53
rect -559 19 -553 53
rect -599 -19 -553 19
rect -599 -53 -593 -19
rect -559 -53 -553 -19
rect -599 -91 -553 -53
rect -599 -125 -593 -91
rect -559 -125 -553 -91
rect -599 -163 -553 -125
rect -599 -197 -593 -163
rect -559 -197 -553 -163
rect -599 -235 -553 -197
rect -599 -269 -593 -235
rect -559 -269 -553 -235
rect -599 -300 -553 -269
rect -503 269 -457 300
rect -503 235 -497 269
rect -463 235 -457 269
rect -503 197 -457 235
rect -503 163 -497 197
rect -463 163 -457 197
rect -503 125 -457 163
rect -503 91 -497 125
rect -463 91 -457 125
rect -503 53 -457 91
rect -503 19 -497 53
rect -463 19 -457 53
rect -503 -19 -457 19
rect -503 -53 -497 -19
rect -463 -53 -457 -19
rect -503 -91 -457 -53
rect -503 -125 -497 -91
rect -463 -125 -457 -91
rect -503 -163 -457 -125
rect -503 -197 -497 -163
rect -463 -197 -457 -163
rect -503 -235 -457 -197
rect -503 -269 -497 -235
rect -463 -269 -457 -235
rect -503 -300 -457 -269
rect -407 269 -361 300
rect -407 235 -401 269
rect -367 235 -361 269
rect -407 197 -361 235
rect -407 163 -401 197
rect -367 163 -361 197
rect -407 125 -361 163
rect -407 91 -401 125
rect -367 91 -361 125
rect -407 53 -361 91
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -91 -361 -53
rect -407 -125 -401 -91
rect -367 -125 -361 -91
rect -407 -163 -361 -125
rect -407 -197 -401 -163
rect -367 -197 -361 -163
rect -407 -235 -361 -197
rect -407 -269 -401 -235
rect -367 -269 -361 -235
rect -407 -300 -361 -269
rect -311 269 -265 300
rect -311 235 -305 269
rect -271 235 -265 269
rect -311 197 -265 235
rect -311 163 -305 197
rect -271 163 -265 197
rect -311 125 -265 163
rect -311 91 -305 125
rect -271 91 -265 125
rect -311 53 -265 91
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -91 -265 -53
rect -311 -125 -305 -91
rect -271 -125 -265 -91
rect -311 -163 -265 -125
rect -311 -197 -305 -163
rect -271 -197 -265 -163
rect -311 -235 -265 -197
rect -311 -269 -305 -235
rect -271 -269 -265 -235
rect -311 -300 -265 -269
rect -215 269 -169 300
rect -215 235 -209 269
rect -175 235 -169 269
rect -215 197 -169 235
rect -215 163 -209 197
rect -175 163 -169 197
rect -215 125 -169 163
rect -215 91 -209 125
rect -175 91 -169 125
rect -215 53 -169 91
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -91 -169 -53
rect -215 -125 -209 -91
rect -175 -125 -169 -91
rect -215 -163 -169 -125
rect -215 -197 -209 -163
rect -175 -197 -169 -163
rect -215 -235 -169 -197
rect -215 -269 -209 -235
rect -175 -269 -169 -235
rect -215 -300 -169 -269
rect -119 269 -73 300
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -300 -73 -269
rect -23 269 23 300
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -300 23 -269
rect 73 269 119 300
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -300 119 -269
rect 169 269 215 300
rect 169 235 175 269
rect 209 235 215 269
rect 169 197 215 235
rect 169 163 175 197
rect 209 163 215 197
rect 169 125 215 163
rect 169 91 175 125
rect 209 91 215 125
rect 169 53 215 91
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -91 215 -53
rect 169 -125 175 -91
rect 209 -125 215 -91
rect 169 -163 215 -125
rect 169 -197 175 -163
rect 209 -197 215 -163
rect 169 -235 215 -197
rect 169 -269 175 -235
rect 209 -269 215 -235
rect 169 -300 215 -269
rect 265 269 311 300
rect 265 235 271 269
rect 305 235 311 269
rect 265 197 311 235
rect 265 163 271 197
rect 305 163 311 197
rect 265 125 311 163
rect 265 91 271 125
rect 305 91 311 125
rect 265 53 311 91
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -91 311 -53
rect 265 -125 271 -91
rect 305 -125 311 -91
rect 265 -163 311 -125
rect 265 -197 271 -163
rect 305 -197 311 -163
rect 265 -235 311 -197
rect 265 -269 271 -235
rect 305 -269 311 -235
rect 265 -300 311 -269
rect 361 269 407 300
rect 361 235 367 269
rect 401 235 407 269
rect 361 197 407 235
rect 361 163 367 197
rect 401 163 407 197
rect 361 125 407 163
rect 361 91 367 125
rect 401 91 407 125
rect 361 53 407 91
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -91 407 -53
rect 361 -125 367 -91
rect 401 -125 407 -91
rect 361 -163 407 -125
rect 361 -197 367 -163
rect 401 -197 407 -163
rect 361 -235 407 -197
rect 361 -269 367 -235
rect 401 -269 407 -235
rect 361 -300 407 -269
rect 457 269 503 300
rect 457 235 463 269
rect 497 235 503 269
rect 457 197 503 235
rect 457 163 463 197
rect 497 163 503 197
rect 457 125 503 163
rect 457 91 463 125
rect 497 91 503 125
rect 457 53 503 91
rect 457 19 463 53
rect 497 19 503 53
rect 457 -19 503 19
rect 457 -53 463 -19
rect 497 -53 503 -19
rect 457 -91 503 -53
rect 457 -125 463 -91
rect 497 -125 503 -91
rect 457 -163 503 -125
rect 457 -197 463 -163
rect 497 -197 503 -163
rect 457 -235 503 -197
rect 457 -269 463 -235
rect 497 -269 503 -235
rect 457 -300 503 -269
rect 553 269 599 300
rect 553 235 559 269
rect 593 235 599 269
rect 553 197 599 235
rect 553 163 559 197
rect 593 163 599 197
rect 553 125 599 163
rect 553 91 559 125
rect 593 91 599 125
rect 553 53 599 91
rect 553 19 559 53
rect 593 19 599 53
rect 553 -19 599 19
rect 553 -53 559 -19
rect 593 -53 599 -19
rect 553 -91 599 -53
rect 553 -125 559 -91
rect 593 -125 599 -91
rect 553 -163 599 -125
rect 553 -197 559 -163
rect 593 -197 599 -163
rect 553 -235 599 -197
rect 553 -269 559 -235
rect 593 -269 599 -235
rect 553 -300 599 -269
rect 649 269 695 300
rect 649 235 655 269
rect 689 235 695 269
rect 649 197 695 235
rect 649 163 655 197
rect 689 163 695 197
rect 649 125 695 163
rect 649 91 655 125
rect 689 91 695 125
rect 649 53 695 91
rect 649 19 655 53
rect 689 19 695 53
rect 649 -19 695 19
rect 649 -53 655 -19
rect 689 -53 695 -19
rect 649 -91 695 -53
rect 649 -125 655 -91
rect 689 -125 695 -91
rect 649 -163 695 -125
rect 649 -197 655 -163
rect 689 -197 695 -163
rect 649 -235 695 -197
rect 649 -269 655 -235
rect 689 -269 695 -235
rect 649 -300 695 -269
rect 745 269 791 300
rect 745 235 751 269
rect 785 235 791 269
rect 745 197 791 235
rect 745 163 751 197
rect 785 163 791 197
rect 745 125 791 163
rect 745 91 751 125
rect 785 91 791 125
rect 745 53 791 91
rect 745 19 751 53
rect 785 19 791 53
rect 745 -19 791 19
rect 745 -53 751 -19
rect 785 -53 791 -19
rect 745 -91 791 -53
rect 745 -125 751 -91
rect 785 -125 791 -91
rect 745 -163 791 -125
rect 745 -197 751 -163
rect 785 -197 791 -163
rect 745 -235 791 -197
rect 745 -269 751 -235
rect 785 -269 791 -235
rect 745 -300 791 -269
rect 841 269 887 300
rect 841 235 847 269
rect 881 235 887 269
rect 841 197 887 235
rect 841 163 847 197
rect 881 163 887 197
rect 841 125 887 163
rect 841 91 847 125
rect 881 91 887 125
rect 841 53 887 91
rect 841 19 847 53
rect 881 19 887 53
rect 841 -19 887 19
rect 841 -53 847 -19
rect 881 -53 887 -19
rect 841 -91 887 -53
rect 841 -125 847 -91
rect 881 -125 887 -91
rect 841 -163 887 -125
rect 841 -197 847 -163
rect 881 -197 887 -163
rect 841 -235 887 -197
rect 841 -269 847 -235
rect 881 -269 887 -235
rect 841 -300 887 -269
rect 937 269 983 300
rect 937 235 943 269
rect 977 235 983 269
rect 937 197 983 235
rect 937 163 943 197
rect 977 163 983 197
rect 937 125 983 163
rect 937 91 943 125
rect 977 91 983 125
rect 937 53 983 91
rect 937 19 943 53
rect 977 19 983 53
rect 937 -19 983 19
rect 937 -53 943 -19
rect 977 -53 983 -19
rect 937 -91 983 -53
rect 937 -125 943 -91
rect 977 -125 983 -91
rect 937 -163 983 -125
rect 937 -197 943 -163
rect 977 -197 983 -163
rect 937 -235 983 -197
rect 937 -269 943 -235
rect 977 -269 983 -235
rect 937 -300 983 -269
rect 1033 269 1079 300
rect 1033 235 1039 269
rect 1073 235 1079 269
rect 1033 197 1079 235
rect 1033 163 1039 197
rect 1073 163 1079 197
rect 1033 125 1079 163
rect 1033 91 1039 125
rect 1073 91 1079 125
rect 1033 53 1079 91
rect 1033 19 1039 53
rect 1073 19 1079 53
rect 1033 -19 1079 19
rect 1033 -53 1039 -19
rect 1073 -53 1079 -19
rect 1033 -91 1079 -53
rect 1033 -125 1039 -91
rect 1073 -125 1079 -91
rect 1033 -163 1079 -125
rect 1033 -197 1039 -163
rect 1073 -197 1079 -163
rect 1033 -235 1079 -197
rect 1033 -269 1039 -235
rect 1073 -269 1079 -235
rect 1033 -300 1079 -269
rect 1129 269 1175 300
rect 1129 235 1135 269
rect 1169 235 1175 269
rect 1129 197 1175 235
rect 1129 163 1135 197
rect 1169 163 1175 197
rect 1129 125 1175 163
rect 1129 91 1135 125
rect 1169 91 1175 125
rect 1129 53 1175 91
rect 1129 19 1135 53
rect 1169 19 1175 53
rect 1129 -19 1175 19
rect 1129 -53 1135 -19
rect 1169 -53 1175 -19
rect 1129 -91 1175 -53
rect 1129 -125 1135 -91
rect 1169 -125 1175 -91
rect 1129 -163 1175 -125
rect 1129 -197 1135 -163
rect 1169 -197 1175 -163
rect 1129 -235 1175 -197
rect 1129 -269 1135 -235
rect 1169 -269 1175 -235
rect 1129 -300 1175 -269
rect 1225 269 1271 300
rect 1225 235 1231 269
rect 1265 235 1271 269
rect 1225 197 1271 235
rect 1225 163 1231 197
rect 1265 163 1271 197
rect 1225 125 1271 163
rect 1225 91 1231 125
rect 1265 91 1271 125
rect 1225 53 1271 91
rect 1225 19 1231 53
rect 1265 19 1271 53
rect 1225 -19 1271 19
rect 1225 -53 1231 -19
rect 1265 -53 1271 -19
rect 1225 -91 1271 -53
rect 1225 -125 1231 -91
rect 1265 -125 1271 -91
rect 1225 -163 1271 -125
rect 1225 -197 1231 -163
rect 1265 -197 1271 -163
rect 1225 -235 1271 -197
rect 1225 -269 1231 -235
rect 1265 -269 1271 -235
rect 1225 -300 1271 -269
rect 1321 269 1367 300
rect 1321 235 1327 269
rect 1361 235 1367 269
rect 1321 197 1367 235
rect 1321 163 1327 197
rect 1361 163 1367 197
rect 1321 125 1367 163
rect 1321 91 1327 125
rect 1361 91 1367 125
rect 1321 53 1367 91
rect 1321 19 1327 53
rect 1361 19 1367 53
rect 1321 -19 1367 19
rect 1321 -53 1327 -19
rect 1361 -53 1367 -19
rect 1321 -91 1367 -53
rect 1321 -125 1327 -91
rect 1361 -125 1367 -91
rect 1321 -163 1367 -125
rect 1321 -197 1327 -163
rect 1361 -197 1367 -163
rect 1321 -235 1367 -197
rect 1321 -269 1327 -235
rect 1361 -269 1367 -235
rect 1321 -300 1367 -269
rect 1417 269 1463 300
rect 1417 235 1423 269
rect 1457 235 1463 269
rect 1417 197 1463 235
rect 1417 163 1423 197
rect 1457 163 1463 197
rect 1417 125 1463 163
rect 1417 91 1423 125
rect 1457 91 1463 125
rect 1417 53 1463 91
rect 1417 19 1423 53
rect 1457 19 1463 53
rect 1417 -19 1463 19
rect 1417 -53 1423 -19
rect 1457 -53 1463 -19
rect 1417 -91 1463 -53
rect 1417 -125 1423 -91
rect 1457 -125 1463 -91
rect 1417 -163 1463 -125
rect 1417 -197 1423 -163
rect 1457 -197 1463 -163
rect 1417 -235 1463 -197
rect 1417 -269 1423 -235
rect 1457 -269 1463 -235
rect 1417 -300 1463 -269
rect 1513 269 1559 300
rect 1513 235 1519 269
rect 1553 235 1559 269
rect 1513 197 1559 235
rect 1513 163 1519 197
rect 1553 163 1559 197
rect 1513 125 1559 163
rect 1513 91 1519 125
rect 1553 91 1559 125
rect 1513 53 1559 91
rect 1513 19 1519 53
rect 1553 19 1559 53
rect 1513 -19 1559 19
rect 1513 -53 1519 -19
rect 1553 -53 1559 -19
rect 1513 -91 1559 -53
rect 1513 -125 1519 -91
rect 1553 -125 1559 -91
rect 1513 -163 1559 -125
rect 1513 -197 1519 -163
rect 1553 -197 1559 -163
rect 1513 -235 1559 -197
rect 1513 -269 1519 -235
rect 1553 -269 1559 -235
rect 1513 -300 1559 -269
rect 1609 269 1655 300
rect 1609 235 1615 269
rect 1649 235 1655 269
rect 1609 197 1655 235
rect 1609 163 1615 197
rect 1649 163 1655 197
rect 1609 125 1655 163
rect 1609 91 1615 125
rect 1649 91 1655 125
rect 1609 53 1655 91
rect 1609 19 1615 53
rect 1649 19 1655 53
rect 1609 -19 1655 19
rect 1609 -53 1615 -19
rect 1649 -53 1655 -19
rect 1609 -91 1655 -53
rect 1609 -125 1615 -91
rect 1649 -125 1655 -91
rect 1609 -163 1655 -125
rect 1609 -197 1615 -163
rect 1649 -197 1655 -163
rect 1609 -235 1655 -197
rect 1609 -269 1615 -235
rect 1649 -269 1655 -235
rect 1609 -300 1655 -269
rect 1705 269 1751 300
rect 1705 235 1711 269
rect 1745 235 1751 269
rect 1705 197 1751 235
rect 1705 163 1711 197
rect 1745 163 1751 197
rect 1705 125 1751 163
rect 1705 91 1711 125
rect 1745 91 1751 125
rect 1705 53 1751 91
rect 1705 19 1711 53
rect 1745 19 1751 53
rect 1705 -19 1751 19
rect 1705 -53 1711 -19
rect 1745 -53 1751 -19
rect 1705 -91 1751 -53
rect 1705 -125 1711 -91
rect 1745 -125 1751 -91
rect 1705 -163 1751 -125
rect 1705 -197 1711 -163
rect 1745 -197 1751 -163
rect 1705 -235 1751 -197
rect 1705 -269 1711 -235
rect 1745 -269 1751 -235
rect 1705 -300 1751 -269
rect 1801 269 1847 300
rect 1801 235 1807 269
rect 1841 235 1847 269
rect 1801 197 1847 235
rect 1801 163 1807 197
rect 1841 163 1847 197
rect 1801 125 1847 163
rect 1801 91 1807 125
rect 1841 91 1847 125
rect 1801 53 1847 91
rect 1801 19 1807 53
rect 1841 19 1847 53
rect 1801 -19 1847 19
rect 1801 -53 1807 -19
rect 1841 -53 1847 -19
rect 1801 -91 1847 -53
rect 1801 -125 1807 -91
rect 1841 -125 1847 -91
rect 1801 -163 1847 -125
rect 1801 -197 1807 -163
rect 1841 -197 1847 -163
rect 1801 -235 1847 -197
rect 1801 -269 1807 -235
rect 1841 -269 1847 -235
rect 1801 -300 1847 -269
rect 1897 269 1943 300
rect 1897 235 1903 269
rect 1937 235 1943 269
rect 1897 197 1943 235
rect 1897 163 1903 197
rect 1937 163 1943 197
rect 1897 125 1943 163
rect 1897 91 1903 125
rect 1937 91 1943 125
rect 1897 53 1943 91
rect 1897 19 1903 53
rect 1937 19 1943 53
rect 1897 -19 1943 19
rect 1897 -53 1903 -19
rect 1937 -53 1943 -19
rect 1897 -91 1943 -53
rect 1897 -125 1903 -91
rect 1937 -125 1943 -91
rect 1897 -163 1943 -125
rect 1897 -197 1903 -163
rect 1937 -197 1943 -163
rect 1897 -235 1943 -197
rect 1897 -269 1903 -235
rect 1937 -269 1943 -235
rect 1897 -300 1943 -269
rect 1993 269 2039 300
rect 1993 235 1999 269
rect 2033 235 2039 269
rect 1993 197 2039 235
rect 1993 163 1999 197
rect 2033 163 2039 197
rect 1993 125 2039 163
rect 1993 91 1999 125
rect 2033 91 2039 125
rect 1993 53 2039 91
rect 1993 19 1999 53
rect 2033 19 2039 53
rect 1993 -19 2039 19
rect 1993 -53 1999 -19
rect 2033 -53 2039 -19
rect 1993 -91 2039 -53
rect 1993 -125 1999 -91
rect 2033 -125 2039 -91
rect 1993 -163 2039 -125
rect 1993 -197 1999 -163
rect 2033 -197 2039 -163
rect 1993 -235 2039 -197
rect 1993 -269 1999 -235
rect 2033 -269 2039 -235
rect 1993 -300 2039 -269
rect -1997 -347 -1939 -341
rect -1997 -381 -1985 -347
rect -1951 -381 -1939 -347
rect -1997 -387 -1939 -381
rect -1805 -347 -1747 -341
rect -1805 -381 -1793 -347
rect -1759 -381 -1747 -347
rect -1805 -387 -1747 -381
rect -1613 -347 -1555 -341
rect -1613 -381 -1601 -347
rect -1567 -381 -1555 -347
rect -1613 -387 -1555 -381
rect -1421 -347 -1363 -341
rect -1421 -381 -1409 -347
rect -1375 -381 -1363 -347
rect -1421 -387 -1363 -381
rect -1229 -347 -1171 -341
rect -1229 -381 -1217 -347
rect -1183 -381 -1171 -347
rect -1229 -387 -1171 -381
rect -1037 -347 -979 -341
rect -1037 -381 -1025 -347
rect -991 -381 -979 -347
rect -1037 -387 -979 -381
rect -845 -347 -787 -341
rect -845 -381 -833 -347
rect -799 -381 -787 -347
rect -845 -387 -787 -381
rect -653 -347 -595 -341
rect -653 -381 -641 -347
rect -607 -381 -595 -347
rect -653 -387 -595 -381
rect -461 -347 -403 -341
rect -461 -381 -449 -347
rect -415 -381 -403 -347
rect -461 -387 -403 -381
rect -269 -347 -211 -341
rect -269 -381 -257 -347
rect -223 -381 -211 -347
rect -269 -387 -211 -381
rect -77 -347 -19 -341
rect -77 -381 -65 -347
rect -31 -381 -19 -347
rect -77 -387 -19 -381
rect 115 -347 173 -341
rect 115 -381 127 -347
rect 161 -381 173 -347
rect 115 -387 173 -381
rect 307 -347 365 -341
rect 307 -381 319 -347
rect 353 -381 365 -347
rect 307 -387 365 -381
rect 499 -347 557 -341
rect 499 -381 511 -347
rect 545 -381 557 -347
rect 499 -387 557 -381
rect 691 -347 749 -341
rect 691 -381 703 -347
rect 737 -381 749 -347
rect 691 -387 749 -381
rect 883 -347 941 -341
rect 883 -381 895 -347
rect 929 -381 941 -347
rect 883 -387 941 -381
rect 1075 -347 1133 -341
rect 1075 -381 1087 -347
rect 1121 -381 1133 -347
rect 1075 -387 1133 -381
rect 1267 -347 1325 -341
rect 1267 -381 1279 -347
rect 1313 -381 1325 -347
rect 1267 -387 1325 -381
rect 1459 -347 1517 -341
rect 1459 -381 1471 -347
rect 1505 -381 1517 -347
rect 1459 -387 1517 -381
rect 1651 -347 1709 -341
rect 1651 -381 1663 -347
rect 1697 -381 1709 -347
rect 1651 -387 1709 -381
rect 1843 -347 1901 -341
rect 1843 -381 1855 -347
rect 1889 -381 1901 -347
rect 1843 -387 1901 -381
<< end >>
