magic
tech sky130A
magscale 1 2
timestamp 1627036492
<< dnwell >>
rect -471 -3014 471 3014
<< nwell >>
rect -551 2808 551 3094
rect -551 -2808 -265 2808
rect 265 -2808 551 2808
rect -551 -3094 551 -2808
<< pwell >>
rect -265 2650 265 2808
rect -265 -2808 265 -2650
<< rpw >>
rect -265 -2650 265 2650
<< psubdiff >>
rect -225 2650 -201 2756
rect 201 2650 225 2756
rect -225 -2756 -201 -2650
rect 201 -2756 225 -2650
<< nsubdiff >>
rect -425 2934 -329 2968
rect 329 2934 425 2968
rect -425 2872 -391 2934
rect 391 2872 425 2934
rect -425 -2934 -391 -2872
rect 391 -2934 425 -2872
rect -425 -2968 -329 -2934
rect 329 -2968 425 -2934
<< psubdiffcont >>
rect -201 2650 201 2756
rect -201 -2756 201 -2650
<< nsubdiffcont >>
rect -329 2934 329 2968
rect -425 -2872 -391 2872
rect 391 -2872 425 2872
rect -329 -2968 329 -2934
<< locali >>
rect -425 2934 -329 2968
rect 329 2934 425 2968
rect -425 2872 -391 2934
rect 391 2872 425 2934
rect -217 2720 -201 2756
rect 201 2720 217 2756
rect -217 2667 -213 2720
rect 213 2667 217 2720
rect -217 2650 -201 2667
rect 201 2650 217 2667
rect -217 -2667 -201 -2650
rect 201 -2667 217 -2650
rect -217 -2720 -213 -2667
rect 213 -2720 217 -2667
rect -217 -2756 -201 -2720
rect 201 -2756 217 -2720
rect -425 -2934 -391 -2872
rect 391 -2934 425 -2872
rect -425 -2968 -329 -2934
rect 329 -2968 425 -2934
<< viali >>
rect -213 2667 -201 2720
rect -201 2667 201 2720
rect 201 2667 213 2720
rect -213 -2720 -201 -2667
rect -201 -2720 201 -2667
rect 201 -2720 213 -2667
<< metal1 >>
rect -225 2720 225 2726
rect -225 2667 -213 2720
rect 213 2667 225 2720
rect -225 2661 225 2667
rect -225 -2667 225 -2661
rect -225 -2720 -213 -2667
rect 213 -2720 225 -2667
rect -225 -2726 225 -2720
<< properties >>
string gencell sky130_fd_pr__res_iso_pw
string FIXED_BBOX -408 -2951 408 2951
string parameters w 2.650 l 26.50 m 1 nx 1 wmin 2.650 lmin 26.50 rho 975 val 10.766k dummy 0 dw 0.25 term 1.0 guard 1 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
