magic
tech sky130A
magscale 1 2
timestamp 1628066849
<< error_p >>
rect 19 492 77 498
rect 19 458 31 492
rect 19 452 77 458
rect -77 -458 -19 -452
rect -77 -492 -65 -458
rect -77 -498 -19 -492
<< pwell >>
rect -263 -630 263 630
<< nmos >>
rect -63 -420 -33 420
rect 33 -420 63 420
<< ndiff >>
rect -125 408 -63 420
rect -125 -408 -113 408
rect -79 -408 -63 408
rect -125 -420 -63 -408
rect -33 408 33 420
rect -33 -408 -17 408
rect 17 -408 33 408
rect -33 -420 33 -408
rect 63 408 125 420
rect 63 -408 79 408
rect 113 -408 125 408
rect 63 -420 125 -408
<< ndiffc >>
rect -113 -408 -79 408
rect -17 -408 17 408
rect 79 -408 113 408
<< psubdiff >>
rect -227 560 -131 594
rect 131 560 227 594
rect -227 498 -193 560
rect 193 498 227 560
rect -227 -560 -193 -498
rect 193 -560 227 -498
rect -227 -594 -131 -560
rect 131 -594 227 -560
<< psubdiffcont >>
rect -131 560 131 594
rect -227 -498 -193 498
rect 193 -498 227 498
rect -131 -594 131 -560
<< poly >>
rect 15 492 81 508
rect 15 458 31 492
rect 65 458 81 492
rect -63 420 -33 446
rect 15 442 81 458
rect 33 420 63 442
rect -63 -442 -33 -420
rect -81 -458 -15 -442
rect 33 -446 63 -420
rect -81 -492 -65 -458
rect -31 -492 -15 -458
rect -81 -508 -15 -492
<< polycont >>
rect 31 458 65 492
rect -65 -492 -31 -458
<< locali >>
rect -227 560 -131 594
rect 131 560 227 594
rect -227 498 -193 560
rect 193 498 227 560
rect 15 458 31 492
rect 65 458 81 492
rect -113 408 -79 424
rect -113 -424 -79 -408
rect -17 408 17 424
rect -17 -424 17 -408
rect 79 408 113 424
rect 79 -424 113 -408
rect -81 -492 -65 -458
rect -31 -492 -15 -458
rect -227 -560 -193 -498
rect 193 -560 227 -498
rect -227 -594 -131 -560
rect 131 -594 227 -560
<< viali >>
rect 31 458 65 492
rect -113 -408 -79 408
rect -17 -408 17 408
rect 79 -408 113 408
rect -65 -492 -31 -458
<< metal1 >>
rect 19 492 77 498
rect 19 458 31 492
rect 65 458 77 492
rect 19 452 77 458
rect -119 408 -73 420
rect -119 -408 -113 408
rect -79 -408 -73 408
rect -119 -420 -73 -408
rect -23 408 23 420
rect -23 -408 -17 408
rect 17 -408 23 408
rect -23 -420 23 -408
rect 73 408 119 420
rect 73 -408 79 408
rect 113 -408 119 408
rect 73 -420 119 -408
rect -77 -458 -19 -452
rect -77 -492 -65 -458
rect -31 -492 -19 -458
rect -77 -498 -19 -492
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -210 -577 210 577
string parameters w 4.2 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
