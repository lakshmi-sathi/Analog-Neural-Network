magic
tech sky130A
magscale 1 2
timestamp 1626798771
<< error_p >>
rect 19 8741 77 8747
rect 19 8707 31 8741
rect 19 8701 77 8707
rect -77 8013 -19 8019
rect -77 7979 -65 8013
rect -77 7973 -19 7979
rect -77 7905 -19 7911
rect -77 7871 -65 7905
rect -77 7865 -19 7871
rect 19 7177 77 7183
rect 19 7143 31 7177
rect 19 7137 77 7143
rect 19 7069 77 7075
rect 19 7035 31 7069
rect 19 7029 77 7035
rect -77 6341 -19 6347
rect -77 6307 -65 6341
rect -77 6301 -19 6307
rect -77 6233 -19 6239
rect -77 6199 -65 6233
rect -77 6193 -19 6199
rect 19 5505 77 5511
rect 19 5471 31 5505
rect 19 5465 77 5471
rect 19 5397 77 5403
rect 19 5363 31 5397
rect 19 5357 77 5363
rect -77 4669 -19 4675
rect -77 4635 -65 4669
rect -77 4629 -19 4635
rect -77 4561 -19 4567
rect -77 4527 -65 4561
rect -77 4521 -19 4527
rect 19 3833 77 3839
rect 19 3799 31 3833
rect 19 3793 77 3799
rect 19 3725 77 3731
rect 19 3691 31 3725
rect 19 3685 77 3691
rect -77 2997 -19 3003
rect -77 2963 -65 2997
rect -77 2957 -19 2963
rect -77 2889 -19 2895
rect -77 2855 -65 2889
rect -77 2849 -19 2855
rect 19 2161 77 2167
rect 19 2127 31 2161
rect 19 2121 77 2127
rect 19 2053 77 2059
rect 19 2019 31 2053
rect 19 2013 77 2019
rect -77 1325 -19 1331
rect -77 1291 -65 1325
rect -77 1285 -19 1291
rect -77 1217 -19 1223
rect -77 1183 -65 1217
rect -77 1177 -19 1183
rect 19 489 77 495
rect 19 455 31 489
rect 19 449 77 455
rect 19 381 77 387
rect 19 347 31 381
rect 19 341 77 347
rect -77 -347 -19 -341
rect -77 -381 -65 -347
rect -77 -387 -19 -381
rect -77 -455 -19 -449
rect -77 -489 -65 -455
rect -77 -495 -19 -489
rect 19 -1183 77 -1177
rect 19 -1217 31 -1183
rect 19 -1223 77 -1217
rect 19 -1291 77 -1285
rect 19 -1325 31 -1291
rect 19 -1331 77 -1325
rect -77 -2019 -19 -2013
rect -77 -2053 -65 -2019
rect -77 -2059 -19 -2053
rect -77 -2127 -19 -2121
rect -77 -2161 -65 -2127
rect -77 -2167 -19 -2161
rect 19 -2855 77 -2849
rect 19 -2889 31 -2855
rect 19 -2895 77 -2889
rect 19 -2963 77 -2957
rect 19 -2997 31 -2963
rect 19 -3003 77 -2997
rect -77 -3691 -19 -3685
rect -77 -3725 -65 -3691
rect -77 -3731 -19 -3725
rect -77 -3799 -19 -3793
rect -77 -3833 -65 -3799
rect -77 -3839 -19 -3833
rect 19 -4527 77 -4521
rect 19 -4561 31 -4527
rect 19 -4567 77 -4561
rect 19 -4635 77 -4629
rect 19 -4669 31 -4635
rect 19 -4675 77 -4669
rect -77 -5363 -19 -5357
rect -77 -5397 -65 -5363
rect -77 -5403 -19 -5397
rect -77 -5471 -19 -5465
rect -77 -5505 -65 -5471
rect -77 -5511 -19 -5505
rect 19 -6199 77 -6193
rect 19 -6233 31 -6199
rect 19 -6239 77 -6233
rect 19 -6307 77 -6301
rect 19 -6341 31 -6307
rect 19 -6347 77 -6341
rect -77 -7035 -19 -7029
rect -77 -7069 -65 -7035
rect -77 -7075 -19 -7069
rect -77 -7143 -19 -7137
rect -77 -7177 -65 -7143
rect -77 -7183 -19 -7177
rect 19 -7871 77 -7865
rect 19 -7905 31 -7871
rect 19 -7911 77 -7905
rect 19 -7979 77 -7973
rect 19 -8013 31 -7979
rect 19 -8019 77 -8013
rect -77 -8707 -19 -8701
rect -77 -8741 -65 -8707
rect -77 -8747 -19 -8741
<< nwell >>
rect -263 -8879 263 8879
<< pmos >>
rect -63 8060 -33 8660
rect 33 8060 63 8660
rect -63 7224 -33 7824
rect 33 7224 63 7824
rect -63 6388 -33 6988
rect 33 6388 63 6988
rect -63 5552 -33 6152
rect 33 5552 63 6152
rect -63 4716 -33 5316
rect 33 4716 63 5316
rect -63 3880 -33 4480
rect 33 3880 63 4480
rect -63 3044 -33 3644
rect 33 3044 63 3644
rect -63 2208 -33 2808
rect 33 2208 63 2808
rect -63 1372 -33 1972
rect 33 1372 63 1972
rect -63 536 -33 1136
rect 33 536 63 1136
rect -63 -300 -33 300
rect 33 -300 63 300
rect -63 -1136 -33 -536
rect 33 -1136 63 -536
rect -63 -1972 -33 -1372
rect 33 -1972 63 -1372
rect -63 -2808 -33 -2208
rect 33 -2808 63 -2208
rect -63 -3644 -33 -3044
rect 33 -3644 63 -3044
rect -63 -4480 -33 -3880
rect 33 -4480 63 -3880
rect -63 -5316 -33 -4716
rect 33 -5316 63 -4716
rect -63 -6152 -33 -5552
rect 33 -6152 63 -5552
rect -63 -6988 -33 -6388
rect 33 -6988 63 -6388
rect -63 -7824 -33 -7224
rect 33 -7824 63 -7224
rect -63 -8660 -33 -8060
rect 33 -8660 63 -8060
<< pdiff >>
rect -125 8648 -63 8660
rect -125 8072 -113 8648
rect -79 8072 -63 8648
rect -125 8060 -63 8072
rect -33 8648 33 8660
rect -33 8072 -17 8648
rect 17 8072 33 8648
rect -33 8060 33 8072
rect 63 8648 125 8660
rect 63 8072 79 8648
rect 113 8072 125 8648
rect 63 8060 125 8072
rect -125 7812 -63 7824
rect -125 7236 -113 7812
rect -79 7236 -63 7812
rect -125 7224 -63 7236
rect -33 7812 33 7824
rect -33 7236 -17 7812
rect 17 7236 33 7812
rect -33 7224 33 7236
rect 63 7812 125 7824
rect 63 7236 79 7812
rect 113 7236 125 7812
rect 63 7224 125 7236
rect -125 6976 -63 6988
rect -125 6400 -113 6976
rect -79 6400 -63 6976
rect -125 6388 -63 6400
rect -33 6976 33 6988
rect -33 6400 -17 6976
rect 17 6400 33 6976
rect -33 6388 33 6400
rect 63 6976 125 6988
rect 63 6400 79 6976
rect 113 6400 125 6976
rect 63 6388 125 6400
rect -125 6140 -63 6152
rect -125 5564 -113 6140
rect -79 5564 -63 6140
rect -125 5552 -63 5564
rect -33 6140 33 6152
rect -33 5564 -17 6140
rect 17 5564 33 6140
rect -33 5552 33 5564
rect 63 6140 125 6152
rect 63 5564 79 6140
rect 113 5564 125 6140
rect 63 5552 125 5564
rect -125 5304 -63 5316
rect -125 4728 -113 5304
rect -79 4728 -63 5304
rect -125 4716 -63 4728
rect -33 5304 33 5316
rect -33 4728 -17 5304
rect 17 4728 33 5304
rect -33 4716 33 4728
rect 63 5304 125 5316
rect 63 4728 79 5304
rect 113 4728 125 5304
rect 63 4716 125 4728
rect -125 4468 -63 4480
rect -125 3892 -113 4468
rect -79 3892 -63 4468
rect -125 3880 -63 3892
rect -33 4468 33 4480
rect -33 3892 -17 4468
rect 17 3892 33 4468
rect -33 3880 33 3892
rect 63 4468 125 4480
rect 63 3892 79 4468
rect 113 3892 125 4468
rect 63 3880 125 3892
rect -125 3632 -63 3644
rect -125 3056 -113 3632
rect -79 3056 -63 3632
rect -125 3044 -63 3056
rect -33 3632 33 3644
rect -33 3056 -17 3632
rect 17 3056 33 3632
rect -33 3044 33 3056
rect 63 3632 125 3644
rect 63 3056 79 3632
rect 113 3056 125 3632
rect 63 3044 125 3056
rect -125 2796 -63 2808
rect -125 2220 -113 2796
rect -79 2220 -63 2796
rect -125 2208 -63 2220
rect -33 2796 33 2808
rect -33 2220 -17 2796
rect 17 2220 33 2796
rect -33 2208 33 2220
rect 63 2796 125 2808
rect 63 2220 79 2796
rect 113 2220 125 2796
rect 63 2208 125 2220
rect -125 1960 -63 1972
rect -125 1384 -113 1960
rect -79 1384 -63 1960
rect -125 1372 -63 1384
rect -33 1960 33 1972
rect -33 1384 -17 1960
rect 17 1384 33 1960
rect -33 1372 33 1384
rect 63 1960 125 1972
rect 63 1384 79 1960
rect 113 1384 125 1960
rect 63 1372 125 1384
rect -125 1124 -63 1136
rect -125 548 -113 1124
rect -79 548 -63 1124
rect -125 536 -63 548
rect -33 1124 33 1136
rect -33 548 -17 1124
rect 17 548 33 1124
rect -33 536 33 548
rect 63 1124 125 1136
rect 63 548 79 1124
rect 113 548 125 1124
rect 63 536 125 548
rect -125 288 -63 300
rect -125 -288 -113 288
rect -79 -288 -63 288
rect -125 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 125 300
rect 63 -288 79 288
rect 113 -288 125 288
rect 63 -300 125 -288
rect -125 -548 -63 -536
rect -125 -1124 -113 -548
rect -79 -1124 -63 -548
rect -125 -1136 -63 -1124
rect -33 -548 33 -536
rect -33 -1124 -17 -548
rect 17 -1124 33 -548
rect -33 -1136 33 -1124
rect 63 -548 125 -536
rect 63 -1124 79 -548
rect 113 -1124 125 -548
rect 63 -1136 125 -1124
rect -125 -1384 -63 -1372
rect -125 -1960 -113 -1384
rect -79 -1960 -63 -1384
rect -125 -1972 -63 -1960
rect -33 -1384 33 -1372
rect -33 -1960 -17 -1384
rect 17 -1960 33 -1384
rect -33 -1972 33 -1960
rect 63 -1384 125 -1372
rect 63 -1960 79 -1384
rect 113 -1960 125 -1384
rect 63 -1972 125 -1960
rect -125 -2220 -63 -2208
rect -125 -2796 -113 -2220
rect -79 -2796 -63 -2220
rect -125 -2808 -63 -2796
rect -33 -2220 33 -2208
rect -33 -2796 -17 -2220
rect 17 -2796 33 -2220
rect -33 -2808 33 -2796
rect 63 -2220 125 -2208
rect 63 -2796 79 -2220
rect 113 -2796 125 -2220
rect 63 -2808 125 -2796
rect -125 -3056 -63 -3044
rect -125 -3632 -113 -3056
rect -79 -3632 -63 -3056
rect -125 -3644 -63 -3632
rect -33 -3056 33 -3044
rect -33 -3632 -17 -3056
rect 17 -3632 33 -3056
rect -33 -3644 33 -3632
rect 63 -3056 125 -3044
rect 63 -3632 79 -3056
rect 113 -3632 125 -3056
rect 63 -3644 125 -3632
rect -125 -3892 -63 -3880
rect -125 -4468 -113 -3892
rect -79 -4468 -63 -3892
rect -125 -4480 -63 -4468
rect -33 -3892 33 -3880
rect -33 -4468 -17 -3892
rect 17 -4468 33 -3892
rect -33 -4480 33 -4468
rect 63 -3892 125 -3880
rect 63 -4468 79 -3892
rect 113 -4468 125 -3892
rect 63 -4480 125 -4468
rect -125 -4728 -63 -4716
rect -125 -5304 -113 -4728
rect -79 -5304 -63 -4728
rect -125 -5316 -63 -5304
rect -33 -4728 33 -4716
rect -33 -5304 -17 -4728
rect 17 -5304 33 -4728
rect -33 -5316 33 -5304
rect 63 -4728 125 -4716
rect 63 -5304 79 -4728
rect 113 -5304 125 -4728
rect 63 -5316 125 -5304
rect -125 -5564 -63 -5552
rect -125 -6140 -113 -5564
rect -79 -6140 -63 -5564
rect -125 -6152 -63 -6140
rect -33 -5564 33 -5552
rect -33 -6140 -17 -5564
rect 17 -6140 33 -5564
rect -33 -6152 33 -6140
rect 63 -5564 125 -5552
rect 63 -6140 79 -5564
rect 113 -6140 125 -5564
rect 63 -6152 125 -6140
rect -125 -6400 -63 -6388
rect -125 -6976 -113 -6400
rect -79 -6976 -63 -6400
rect -125 -6988 -63 -6976
rect -33 -6400 33 -6388
rect -33 -6976 -17 -6400
rect 17 -6976 33 -6400
rect -33 -6988 33 -6976
rect 63 -6400 125 -6388
rect 63 -6976 79 -6400
rect 113 -6976 125 -6400
rect 63 -6988 125 -6976
rect -125 -7236 -63 -7224
rect -125 -7812 -113 -7236
rect -79 -7812 -63 -7236
rect -125 -7824 -63 -7812
rect -33 -7236 33 -7224
rect -33 -7812 -17 -7236
rect 17 -7812 33 -7236
rect -33 -7824 33 -7812
rect 63 -7236 125 -7224
rect 63 -7812 79 -7236
rect 113 -7812 125 -7236
rect 63 -7824 125 -7812
rect -125 -8072 -63 -8060
rect -125 -8648 -113 -8072
rect -79 -8648 -63 -8072
rect -125 -8660 -63 -8648
rect -33 -8072 33 -8060
rect -33 -8648 -17 -8072
rect 17 -8648 33 -8072
rect -33 -8660 33 -8648
rect 63 -8072 125 -8060
rect 63 -8648 79 -8072
rect 113 -8648 125 -8072
rect 63 -8660 125 -8648
<< pdiffc >>
rect -113 8072 -79 8648
rect -17 8072 17 8648
rect 79 8072 113 8648
rect -113 7236 -79 7812
rect -17 7236 17 7812
rect 79 7236 113 7812
rect -113 6400 -79 6976
rect -17 6400 17 6976
rect 79 6400 113 6976
rect -113 5564 -79 6140
rect -17 5564 17 6140
rect 79 5564 113 6140
rect -113 4728 -79 5304
rect -17 4728 17 5304
rect 79 4728 113 5304
rect -113 3892 -79 4468
rect -17 3892 17 4468
rect 79 3892 113 4468
rect -113 3056 -79 3632
rect -17 3056 17 3632
rect 79 3056 113 3632
rect -113 2220 -79 2796
rect -17 2220 17 2796
rect 79 2220 113 2796
rect -113 1384 -79 1960
rect -17 1384 17 1960
rect 79 1384 113 1960
rect -113 548 -79 1124
rect -17 548 17 1124
rect 79 548 113 1124
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect -113 -1124 -79 -548
rect -17 -1124 17 -548
rect 79 -1124 113 -548
rect -113 -1960 -79 -1384
rect -17 -1960 17 -1384
rect 79 -1960 113 -1384
rect -113 -2796 -79 -2220
rect -17 -2796 17 -2220
rect 79 -2796 113 -2220
rect -113 -3632 -79 -3056
rect -17 -3632 17 -3056
rect 79 -3632 113 -3056
rect -113 -4468 -79 -3892
rect -17 -4468 17 -3892
rect 79 -4468 113 -3892
rect -113 -5304 -79 -4728
rect -17 -5304 17 -4728
rect 79 -5304 113 -4728
rect -113 -6140 -79 -5564
rect -17 -6140 17 -5564
rect 79 -6140 113 -5564
rect -113 -6976 -79 -6400
rect -17 -6976 17 -6400
rect 79 -6976 113 -6400
rect -113 -7812 -79 -7236
rect -17 -7812 17 -7236
rect 79 -7812 113 -7236
rect -113 -8648 -79 -8072
rect -17 -8648 17 -8072
rect 79 -8648 113 -8072
<< nsubdiff >>
rect -227 8809 -131 8843
rect 131 8809 227 8843
rect -227 8747 -193 8809
rect 193 8747 227 8809
rect -227 -8809 -193 -8747
rect 193 -8809 227 -8747
rect -227 -8843 -131 -8809
rect 131 -8843 227 -8809
<< nsubdiffcont >>
rect -131 8809 131 8843
rect -227 -8747 -193 8747
rect 193 -8747 227 8747
rect -131 -8843 131 -8809
<< poly >>
rect 15 8741 81 8757
rect 15 8707 31 8741
rect 65 8707 81 8741
rect 15 8691 81 8707
rect -63 8660 -33 8686
rect 33 8660 63 8691
rect -63 8029 -33 8060
rect 33 8034 63 8060
rect -81 8013 -15 8029
rect -81 7979 -65 8013
rect -31 7979 -15 8013
rect -81 7963 -15 7979
rect -81 7905 -15 7921
rect -81 7871 -65 7905
rect -31 7871 -15 7905
rect -81 7855 -15 7871
rect -63 7824 -33 7855
rect 33 7824 63 7850
rect -63 7198 -33 7224
rect 33 7193 63 7224
rect 15 7177 81 7193
rect 15 7143 31 7177
rect 65 7143 81 7177
rect 15 7127 81 7143
rect 15 7069 81 7085
rect 15 7035 31 7069
rect 65 7035 81 7069
rect 15 7019 81 7035
rect -63 6988 -33 7014
rect 33 6988 63 7019
rect -63 6357 -33 6388
rect 33 6362 63 6388
rect -81 6341 -15 6357
rect -81 6307 -65 6341
rect -31 6307 -15 6341
rect -81 6291 -15 6307
rect -81 6233 -15 6249
rect -81 6199 -65 6233
rect -31 6199 -15 6233
rect -81 6183 -15 6199
rect -63 6152 -33 6183
rect 33 6152 63 6178
rect -63 5526 -33 5552
rect 33 5521 63 5552
rect 15 5505 81 5521
rect 15 5471 31 5505
rect 65 5471 81 5505
rect 15 5455 81 5471
rect 15 5397 81 5413
rect 15 5363 31 5397
rect 65 5363 81 5397
rect 15 5347 81 5363
rect -63 5316 -33 5342
rect 33 5316 63 5347
rect -63 4685 -33 4716
rect 33 4690 63 4716
rect -81 4669 -15 4685
rect -81 4635 -65 4669
rect -31 4635 -15 4669
rect -81 4619 -15 4635
rect -81 4561 -15 4577
rect -81 4527 -65 4561
rect -31 4527 -15 4561
rect -81 4511 -15 4527
rect -63 4480 -33 4511
rect 33 4480 63 4506
rect -63 3854 -33 3880
rect 33 3849 63 3880
rect 15 3833 81 3849
rect 15 3799 31 3833
rect 65 3799 81 3833
rect 15 3783 81 3799
rect 15 3725 81 3741
rect 15 3691 31 3725
rect 65 3691 81 3725
rect 15 3675 81 3691
rect -63 3644 -33 3670
rect 33 3644 63 3675
rect -63 3013 -33 3044
rect 33 3018 63 3044
rect -81 2997 -15 3013
rect -81 2963 -65 2997
rect -31 2963 -15 2997
rect -81 2947 -15 2963
rect -81 2889 -15 2905
rect -81 2855 -65 2889
rect -31 2855 -15 2889
rect -81 2839 -15 2855
rect -63 2808 -33 2839
rect 33 2808 63 2834
rect -63 2182 -33 2208
rect 33 2177 63 2208
rect 15 2161 81 2177
rect 15 2127 31 2161
rect 65 2127 81 2161
rect 15 2111 81 2127
rect 15 2053 81 2069
rect 15 2019 31 2053
rect 65 2019 81 2053
rect 15 2003 81 2019
rect -63 1972 -33 1998
rect 33 1972 63 2003
rect -63 1341 -33 1372
rect 33 1346 63 1372
rect -81 1325 -15 1341
rect -81 1291 -65 1325
rect -31 1291 -15 1325
rect -81 1275 -15 1291
rect -81 1217 -15 1233
rect -81 1183 -65 1217
rect -31 1183 -15 1217
rect -81 1167 -15 1183
rect -63 1136 -33 1167
rect 33 1136 63 1162
rect -63 510 -33 536
rect 33 505 63 536
rect 15 489 81 505
rect 15 455 31 489
rect 65 455 81 489
rect 15 439 81 455
rect 15 381 81 397
rect 15 347 31 381
rect 65 347 81 381
rect 15 331 81 347
rect -63 300 -33 326
rect 33 300 63 331
rect -63 -331 -33 -300
rect 33 -326 63 -300
rect -81 -347 -15 -331
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect -81 -397 -15 -381
rect -81 -455 -15 -439
rect -81 -489 -65 -455
rect -31 -489 -15 -455
rect -81 -505 -15 -489
rect -63 -536 -33 -505
rect 33 -536 63 -510
rect -63 -1162 -33 -1136
rect 33 -1167 63 -1136
rect 15 -1183 81 -1167
rect 15 -1217 31 -1183
rect 65 -1217 81 -1183
rect 15 -1233 81 -1217
rect 15 -1291 81 -1275
rect 15 -1325 31 -1291
rect 65 -1325 81 -1291
rect 15 -1341 81 -1325
rect -63 -1372 -33 -1346
rect 33 -1372 63 -1341
rect -63 -2003 -33 -1972
rect 33 -1998 63 -1972
rect -81 -2019 -15 -2003
rect -81 -2053 -65 -2019
rect -31 -2053 -15 -2019
rect -81 -2069 -15 -2053
rect -81 -2127 -15 -2111
rect -81 -2161 -65 -2127
rect -31 -2161 -15 -2127
rect -81 -2177 -15 -2161
rect -63 -2208 -33 -2177
rect 33 -2208 63 -2182
rect -63 -2834 -33 -2808
rect 33 -2839 63 -2808
rect 15 -2855 81 -2839
rect 15 -2889 31 -2855
rect 65 -2889 81 -2855
rect 15 -2905 81 -2889
rect 15 -2963 81 -2947
rect 15 -2997 31 -2963
rect 65 -2997 81 -2963
rect 15 -3013 81 -2997
rect -63 -3044 -33 -3018
rect 33 -3044 63 -3013
rect -63 -3675 -33 -3644
rect 33 -3670 63 -3644
rect -81 -3691 -15 -3675
rect -81 -3725 -65 -3691
rect -31 -3725 -15 -3691
rect -81 -3741 -15 -3725
rect -81 -3799 -15 -3783
rect -81 -3833 -65 -3799
rect -31 -3833 -15 -3799
rect -81 -3849 -15 -3833
rect -63 -3880 -33 -3849
rect 33 -3880 63 -3854
rect -63 -4506 -33 -4480
rect 33 -4511 63 -4480
rect 15 -4527 81 -4511
rect 15 -4561 31 -4527
rect 65 -4561 81 -4527
rect 15 -4577 81 -4561
rect 15 -4635 81 -4619
rect 15 -4669 31 -4635
rect 65 -4669 81 -4635
rect 15 -4685 81 -4669
rect -63 -4716 -33 -4690
rect 33 -4716 63 -4685
rect -63 -5347 -33 -5316
rect 33 -5342 63 -5316
rect -81 -5363 -15 -5347
rect -81 -5397 -65 -5363
rect -31 -5397 -15 -5363
rect -81 -5413 -15 -5397
rect -81 -5471 -15 -5455
rect -81 -5505 -65 -5471
rect -31 -5505 -15 -5471
rect -81 -5521 -15 -5505
rect -63 -5552 -33 -5521
rect 33 -5552 63 -5526
rect -63 -6178 -33 -6152
rect 33 -6183 63 -6152
rect 15 -6199 81 -6183
rect 15 -6233 31 -6199
rect 65 -6233 81 -6199
rect 15 -6249 81 -6233
rect 15 -6307 81 -6291
rect 15 -6341 31 -6307
rect 65 -6341 81 -6307
rect 15 -6357 81 -6341
rect -63 -6388 -33 -6362
rect 33 -6388 63 -6357
rect -63 -7019 -33 -6988
rect 33 -7014 63 -6988
rect -81 -7035 -15 -7019
rect -81 -7069 -65 -7035
rect -31 -7069 -15 -7035
rect -81 -7085 -15 -7069
rect -81 -7143 -15 -7127
rect -81 -7177 -65 -7143
rect -31 -7177 -15 -7143
rect -81 -7193 -15 -7177
rect -63 -7224 -33 -7193
rect 33 -7224 63 -7198
rect -63 -7850 -33 -7824
rect 33 -7855 63 -7824
rect 15 -7871 81 -7855
rect 15 -7905 31 -7871
rect 65 -7905 81 -7871
rect 15 -7921 81 -7905
rect 15 -7979 81 -7963
rect 15 -8013 31 -7979
rect 65 -8013 81 -7979
rect 15 -8029 81 -8013
rect -63 -8060 -33 -8034
rect 33 -8060 63 -8029
rect -63 -8691 -33 -8660
rect 33 -8686 63 -8660
rect -81 -8707 -15 -8691
rect -81 -8741 -65 -8707
rect -31 -8741 -15 -8707
rect -81 -8757 -15 -8741
<< polycont >>
rect 31 8707 65 8741
rect -65 7979 -31 8013
rect -65 7871 -31 7905
rect 31 7143 65 7177
rect 31 7035 65 7069
rect -65 6307 -31 6341
rect -65 6199 -31 6233
rect 31 5471 65 5505
rect 31 5363 65 5397
rect -65 4635 -31 4669
rect -65 4527 -31 4561
rect 31 3799 65 3833
rect 31 3691 65 3725
rect -65 2963 -31 2997
rect -65 2855 -31 2889
rect 31 2127 65 2161
rect 31 2019 65 2053
rect -65 1291 -31 1325
rect -65 1183 -31 1217
rect 31 455 65 489
rect 31 347 65 381
rect -65 -381 -31 -347
rect -65 -489 -31 -455
rect 31 -1217 65 -1183
rect 31 -1325 65 -1291
rect -65 -2053 -31 -2019
rect -65 -2161 -31 -2127
rect 31 -2889 65 -2855
rect 31 -2997 65 -2963
rect -65 -3725 -31 -3691
rect -65 -3833 -31 -3799
rect 31 -4561 65 -4527
rect 31 -4669 65 -4635
rect -65 -5397 -31 -5363
rect -65 -5505 -31 -5471
rect 31 -6233 65 -6199
rect 31 -6341 65 -6307
rect -65 -7069 -31 -7035
rect -65 -7177 -31 -7143
rect 31 -7905 65 -7871
rect 31 -8013 65 -7979
rect -65 -8741 -31 -8707
<< locali >>
rect -227 8809 -131 8843
rect 131 8809 227 8843
rect -227 8747 -193 8809
rect 193 8747 227 8809
rect 15 8707 31 8741
rect 65 8707 81 8741
rect -113 8648 -79 8664
rect -113 8056 -79 8072
rect -17 8648 17 8664
rect -17 8056 17 8072
rect 79 8648 113 8664
rect 79 8056 113 8072
rect -81 7979 -65 8013
rect -31 7979 -15 8013
rect -81 7871 -65 7905
rect -31 7871 -15 7905
rect -113 7812 -79 7828
rect -113 7220 -79 7236
rect -17 7812 17 7828
rect -17 7220 17 7236
rect 79 7812 113 7828
rect 79 7220 113 7236
rect 15 7143 31 7177
rect 65 7143 81 7177
rect 15 7035 31 7069
rect 65 7035 81 7069
rect -113 6976 -79 6992
rect -113 6384 -79 6400
rect -17 6976 17 6992
rect -17 6384 17 6400
rect 79 6976 113 6992
rect 79 6384 113 6400
rect -81 6307 -65 6341
rect -31 6307 -15 6341
rect -81 6199 -65 6233
rect -31 6199 -15 6233
rect -113 6140 -79 6156
rect -113 5548 -79 5564
rect -17 6140 17 6156
rect -17 5548 17 5564
rect 79 6140 113 6156
rect 79 5548 113 5564
rect 15 5471 31 5505
rect 65 5471 81 5505
rect 15 5363 31 5397
rect 65 5363 81 5397
rect -113 5304 -79 5320
rect -113 4712 -79 4728
rect -17 5304 17 5320
rect -17 4712 17 4728
rect 79 5304 113 5320
rect 79 4712 113 4728
rect -81 4635 -65 4669
rect -31 4635 -15 4669
rect -81 4527 -65 4561
rect -31 4527 -15 4561
rect -113 4468 -79 4484
rect -113 3876 -79 3892
rect -17 4468 17 4484
rect -17 3876 17 3892
rect 79 4468 113 4484
rect 79 3876 113 3892
rect 15 3799 31 3833
rect 65 3799 81 3833
rect 15 3691 31 3725
rect 65 3691 81 3725
rect -113 3632 -79 3648
rect -113 3040 -79 3056
rect -17 3632 17 3648
rect -17 3040 17 3056
rect 79 3632 113 3648
rect 79 3040 113 3056
rect -81 2963 -65 2997
rect -31 2963 -15 2997
rect -81 2855 -65 2889
rect -31 2855 -15 2889
rect -113 2796 -79 2812
rect -113 2204 -79 2220
rect -17 2796 17 2812
rect -17 2204 17 2220
rect 79 2796 113 2812
rect 79 2204 113 2220
rect 15 2127 31 2161
rect 65 2127 81 2161
rect 15 2019 31 2053
rect 65 2019 81 2053
rect -113 1960 -79 1976
rect -113 1368 -79 1384
rect -17 1960 17 1976
rect -17 1368 17 1384
rect 79 1960 113 1976
rect 79 1368 113 1384
rect -81 1291 -65 1325
rect -31 1291 -15 1325
rect -81 1183 -65 1217
rect -31 1183 -15 1217
rect -113 1124 -79 1140
rect -113 532 -79 548
rect -17 1124 17 1140
rect -17 532 17 548
rect 79 1124 113 1140
rect 79 532 113 548
rect 15 455 31 489
rect 65 455 81 489
rect 15 347 31 381
rect 65 347 81 381
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect -81 -489 -65 -455
rect -31 -489 -15 -455
rect -113 -548 -79 -532
rect -113 -1140 -79 -1124
rect -17 -548 17 -532
rect -17 -1140 17 -1124
rect 79 -548 113 -532
rect 79 -1140 113 -1124
rect 15 -1217 31 -1183
rect 65 -1217 81 -1183
rect 15 -1325 31 -1291
rect 65 -1325 81 -1291
rect -113 -1384 -79 -1368
rect -113 -1976 -79 -1960
rect -17 -1384 17 -1368
rect -17 -1976 17 -1960
rect 79 -1384 113 -1368
rect 79 -1976 113 -1960
rect -81 -2053 -65 -2019
rect -31 -2053 -15 -2019
rect -81 -2161 -65 -2127
rect -31 -2161 -15 -2127
rect -113 -2220 -79 -2204
rect -113 -2812 -79 -2796
rect -17 -2220 17 -2204
rect -17 -2812 17 -2796
rect 79 -2220 113 -2204
rect 79 -2812 113 -2796
rect 15 -2889 31 -2855
rect 65 -2889 81 -2855
rect 15 -2997 31 -2963
rect 65 -2997 81 -2963
rect -113 -3056 -79 -3040
rect -113 -3648 -79 -3632
rect -17 -3056 17 -3040
rect -17 -3648 17 -3632
rect 79 -3056 113 -3040
rect 79 -3648 113 -3632
rect -81 -3725 -65 -3691
rect -31 -3725 -15 -3691
rect -81 -3833 -65 -3799
rect -31 -3833 -15 -3799
rect -113 -3892 -79 -3876
rect -113 -4484 -79 -4468
rect -17 -3892 17 -3876
rect -17 -4484 17 -4468
rect 79 -3892 113 -3876
rect 79 -4484 113 -4468
rect 15 -4561 31 -4527
rect 65 -4561 81 -4527
rect 15 -4669 31 -4635
rect 65 -4669 81 -4635
rect -113 -4728 -79 -4712
rect -113 -5320 -79 -5304
rect -17 -4728 17 -4712
rect -17 -5320 17 -5304
rect 79 -4728 113 -4712
rect 79 -5320 113 -5304
rect -81 -5397 -65 -5363
rect -31 -5397 -15 -5363
rect -81 -5505 -65 -5471
rect -31 -5505 -15 -5471
rect -113 -5564 -79 -5548
rect -113 -6156 -79 -6140
rect -17 -5564 17 -5548
rect -17 -6156 17 -6140
rect 79 -5564 113 -5548
rect 79 -6156 113 -6140
rect 15 -6233 31 -6199
rect 65 -6233 81 -6199
rect 15 -6341 31 -6307
rect 65 -6341 81 -6307
rect -113 -6400 -79 -6384
rect -113 -6992 -79 -6976
rect -17 -6400 17 -6384
rect -17 -6992 17 -6976
rect 79 -6400 113 -6384
rect 79 -6992 113 -6976
rect -81 -7069 -65 -7035
rect -31 -7069 -15 -7035
rect -81 -7177 -65 -7143
rect -31 -7177 -15 -7143
rect -113 -7236 -79 -7220
rect -113 -7828 -79 -7812
rect -17 -7236 17 -7220
rect -17 -7828 17 -7812
rect 79 -7236 113 -7220
rect 79 -7828 113 -7812
rect 15 -7905 31 -7871
rect 65 -7905 81 -7871
rect 15 -8013 31 -7979
rect 65 -8013 81 -7979
rect -113 -8072 -79 -8056
rect -113 -8664 -79 -8648
rect -17 -8072 17 -8056
rect -17 -8664 17 -8648
rect 79 -8072 113 -8056
rect 79 -8664 113 -8648
rect -81 -8741 -65 -8707
rect -31 -8741 -15 -8707
rect -227 -8809 -193 -8747
rect 193 -8809 227 -8747
rect -227 -8843 -131 -8809
rect 131 -8843 227 -8809
<< viali >>
rect 31 8707 65 8741
rect -113 8072 -79 8648
rect -17 8072 17 8648
rect 79 8072 113 8648
rect -65 7979 -31 8013
rect -65 7871 -31 7905
rect -113 7236 -79 7812
rect -17 7236 17 7812
rect 79 7236 113 7812
rect 31 7143 65 7177
rect 31 7035 65 7069
rect -113 6400 -79 6976
rect -17 6400 17 6976
rect 79 6400 113 6976
rect -65 6307 -31 6341
rect -65 6199 -31 6233
rect -113 5564 -79 6140
rect -17 5564 17 6140
rect 79 5564 113 6140
rect 31 5471 65 5505
rect 31 5363 65 5397
rect -113 4728 -79 5304
rect -17 4728 17 5304
rect 79 4728 113 5304
rect -65 4635 -31 4669
rect -65 4527 -31 4561
rect -113 3892 -79 4468
rect -17 3892 17 4468
rect 79 3892 113 4468
rect 31 3799 65 3833
rect 31 3691 65 3725
rect -113 3056 -79 3632
rect -17 3056 17 3632
rect 79 3056 113 3632
rect -65 2963 -31 2997
rect -65 2855 -31 2889
rect -113 2220 -79 2796
rect -17 2220 17 2796
rect 79 2220 113 2796
rect 31 2127 65 2161
rect 31 2019 65 2053
rect -113 1384 -79 1960
rect -17 1384 17 1960
rect 79 1384 113 1960
rect -65 1291 -31 1325
rect -65 1183 -31 1217
rect -113 548 -79 1124
rect -17 548 17 1124
rect 79 548 113 1124
rect 31 455 65 489
rect 31 347 65 381
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect -65 -381 -31 -347
rect -65 -489 -31 -455
rect -113 -1124 -79 -548
rect -17 -1124 17 -548
rect 79 -1124 113 -548
rect 31 -1217 65 -1183
rect 31 -1325 65 -1291
rect -113 -1960 -79 -1384
rect -17 -1960 17 -1384
rect 79 -1960 113 -1384
rect -65 -2053 -31 -2019
rect -65 -2161 -31 -2127
rect -113 -2796 -79 -2220
rect -17 -2796 17 -2220
rect 79 -2796 113 -2220
rect 31 -2889 65 -2855
rect 31 -2997 65 -2963
rect -113 -3632 -79 -3056
rect -17 -3632 17 -3056
rect 79 -3632 113 -3056
rect -65 -3725 -31 -3691
rect -65 -3833 -31 -3799
rect -113 -4468 -79 -3892
rect -17 -4468 17 -3892
rect 79 -4468 113 -3892
rect 31 -4561 65 -4527
rect 31 -4669 65 -4635
rect -113 -5304 -79 -4728
rect -17 -5304 17 -4728
rect 79 -5304 113 -4728
rect -65 -5397 -31 -5363
rect -65 -5505 -31 -5471
rect -113 -6140 -79 -5564
rect -17 -6140 17 -5564
rect 79 -6140 113 -5564
rect 31 -6233 65 -6199
rect 31 -6341 65 -6307
rect -113 -6976 -79 -6400
rect -17 -6976 17 -6400
rect 79 -6976 113 -6400
rect -65 -7069 -31 -7035
rect -65 -7177 -31 -7143
rect -113 -7812 -79 -7236
rect -17 -7812 17 -7236
rect 79 -7812 113 -7236
rect 31 -7905 65 -7871
rect 31 -8013 65 -7979
rect -113 -8648 -79 -8072
rect -17 -8648 17 -8072
rect 79 -8648 113 -8072
rect -65 -8741 -31 -8707
<< metal1 >>
rect 19 8741 77 8747
rect 19 8707 31 8741
rect 65 8707 77 8741
rect 19 8701 77 8707
rect -119 8648 -73 8660
rect -119 8072 -113 8648
rect -79 8072 -73 8648
rect -119 8060 -73 8072
rect -23 8648 23 8660
rect -23 8072 -17 8648
rect 17 8072 23 8648
rect -23 8060 23 8072
rect 73 8648 119 8660
rect 73 8072 79 8648
rect 113 8072 119 8648
rect 73 8060 119 8072
rect -77 8013 -19 8019
rect -77 7979 -65 8013
rect -31 7979 -19 8013
rect -77 7973 -19 7979
rect -77 7905 -19 7911
rect -77 7871 -65 7905
rect -31 7871 -19 7905
rect -77 7865 -19 7871
rect -119 7812 -73 7824
rect -119 7236 -113 7812
rect -79 7236 -73 7812
rect -119 7224 -73 7236
rect -23 7812 23 7824
rect -23 7236 -17 7812
rect 17 7236 23 7812
rect -23 7224 23 7236
rect 73 7812 119 7824
rect 73 7236 79 7812
rect 113 7236 119 7812
rect 73 7224 119 7236
rect 19 7177 77 7183
rect 19 7143 31 7177
rect 65 7143 77 7177
rect 19 7137 77 7143
rect 19 7069 77 7075
rect 19 7035 31 7069
rect 65 7035 77 7069
rect 19 7029 77 7035
rect -119 6976 -73 6988
rect -119 6400 -113 6976
rect -79 6400 -73 6976
rect -119 6388 -73 6400
rect -23 6976 23 6988
rect -23 6400 -17 6976
rect 17 6400 23 6976
rect -23 6388 23 6400
rect 73 6976 119 6988
rect 73 6400 79 6976
rect 113 6400 119 6976
rect 73 6388 119 6400
rect -77 6341 -19 6347
rect -77 6307 -65 6341
rect -31 6307 -19 6341
rect -77 6301 -19 6307
rect -77 6233 -19 6239
rect -77 6199 -65 6233
rect -31 6199 -19 6233
rect -77 6193 -19 6199
rect -119 6140 -73 6152
rect -119 5564 -113 6140
rect -79 5564 -73 6140
rect -119 5552 -73 5564
rect -23 6140 23 6152
rect -23 5564 -17 6140
rect 17 5564 23 6140
rect -23 5552 23 5564
rect 73 6140 119 6152
rect 73 5564 79 6140
rect 113 5564 119 6140
rect 73 5552 119 5564
rect 19 5505 77 5511
rect 19 5471 31 5505
rect 65 5471 77 5505
rect 19 5465 77 5471
rect 19 5397 77 5403
rect 19 5363 31 5397
rect 65 5363 77 5397
rect 19 5357 77 5363
rect -119 5304 -73 5316
rect -119 4728 -113 5304
rect -79 4728 -73 5304
rect -119 4716 -73 4728
rect -23 5304 23 5316
rect -23 4728 -17 5304
rect 17 4728 23 5304
rect -23 4716 23 4728
rect 73 5304 119 5316
rect 73 4728 79 5304
rect 113 4728 119 5304
rect 73 4716 119 4728
rect -77 4669 -19 4675
rect -77 4635 -65 4669
rect -31 4635 -19 4669
rect -77 4629 -19 4635
rect -77 4561 -19 4567
rect -77 4527 -65 4561
rect -31 4527 -19 4561
rect -77 4521 -19 4527
rect -119 4468 -73 4480
rect -119 3892 -113 4468
rect -79 3892 -73 4468
rect -119 3880 -73 3892
rect -23 4468 23 4480
rect -23 3892 -17 4468
rect 17 3892 23 4468
rect -23 3880 23 3892
rect 73 4468 119 4480
rect 73 3892 79 4468
rect 113 3892 119 4468
rect 73 3880 119 3892
rect 19 3833 77 3839
rect 19 3799 31 3833
rect 65 3799 77 3833
rect 19 3793 77 3799
rect 19 3725 77 3731
rect 19 3691 31 3725
rect 65 3691 77 3725
rect 19 3685 77 3691
rect -119 3632 -73 3644
rect -119 3056 -113 3632
rect -79 3056 -73 3632
rect -119 3044 -73 3056
rect -23 3632 23 3644
rect -23 3056 -17 3632
rect 17 3056 23 3632
rect -23 3044 23 3056
rect 73 3632 119 3644
rect 73 3056 79 3632
rect 113 3056 119 3632
rect 73 3044 119 3056
rect -77 2997 -19 3003
rect -77 2963 -65 2997
rect -31 2963 -19 2997
rect -77 2957 -19 2963
rect -77 2889 -19 2895
rect -77 2855 -65 2889
rect -31 2855 -19 2889
rect -77 2849 -19 2855
rect -119 2796 -73 2808
rect -119 2220 -113 2796
rect -79 2220 -73 2796
rect -119 2208 -73 2220
rect -23 2796 23 2808
rect -23 2220 -17 2796
rect 17 2220 23 2796
rect -23 2208 23 2220
rect 73 2796 119 2808
rect 73 2220 79 2796
rect 113 2220 119 2796
rect 73 2208 119 2220
rect 19 2161 77 2167
rect 19 2127 31 2161
rect 65 2127 77 2161
rect 19 2121 77 2127
rect 19 2053 77 2059
rect 19 2019 31 2053
rect 65 2019 77 2053
rect 19 2013 77 2019
rect -119 1960 -73 1972
rect -119 1384 -113 1960
rect -79 1384 -73 1960
rect -119 1372 -73 1384
rect -23 1960 23 1972
rect -23 1384 -17 1960
rect 17 1384 23 1960
rect -23 1372 23 1384
rect 73 1960 119 1972
rect 73 1384 79 1960
rect 113 1384 119 1960
rect 73 1372 119 1384
rect -77 1325 -19 1331
rect -77 1291 -65 1325
rect -31 1291 -19 1325
rect -77 1285 -19 1291
rect -77 1217 -19 1223
rect -77 1183 -65 1217
rect -31 1183 -19 1217
rect -77 1177 -19 1183
rect -119 1124 -73 1136
rect -119 548 -113 1124
rect -79 548 -73 1124
rect -119 536 -73 548
rect -23 1124 23 1136
rect -23 548 -17 1124
rect 17 548 23 1124
rect -23 536 23 548
rect 73 1124 119 1136
rect 73 548 79 1124
rect 113 548 119 1124
rect 73 536 119 548
rect 19 489 77 495
rect 19 455 31 489
rect 65 455 77 489
rect 19 449 77 455
rect 19 381 77 387
rect 19 347 31 381
rect 65 347 77 381
rect 19 341 77 347
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect -77 -347 -19 -341
rect -77 -381 -65 -347
rect -31 -381 -19 -347
rect -77 -387 -19 -381
rect -77 -455 -19 -449
rect -77 -489 -65 -455
rect -31 -489 -19 -455
rect -77 -495 -19 -489
rect -119 -548 -73 -536
rect -119 -1124 -113 -548
rect -79 -1124 -73 -548
rect -119 -1136 -73 -1124
rect -23 -548 23 -536
rect -23 -1124 -17 -548
rect 17 -1124 23 -548
rect -23 -1136 23 -1124
rect 73 -548 119 -536
rect 73 -1124 79 -548
rect 113 -1124 119 -548
rect 73 -1136 119 -1124
rect 19 -1183 77 -1177
rect 19 -1217 31 -1183
rect 65 -1217 77 -1183
rect 19 -1223 77 -1217
rect 19 -1291 77 -1285
rect 19 -1325 31 -1291
rect 65 -1325 77 -1291
rect 19 -1331 77 -1325
rect -119 -1384 -73 -1372
rect -119 -1960 -113 -1384
rect -79 -1960 -73 -1384
rect -119 -1972 -73 -1960
rect -23 -1384 23 -1372
rect -23 -1960 -17 -1384
rect 17 -1960 23 -1384
rect -23 -1972 23 -1960
rect 73 -1384 119 -1372
rect 73 -1960 79 -1384
rect 113 -1960 119 -1384
rect 73 -1972 119 -1960
rect -77 -2019 -19 -2013
rect -77 -2053 -65 -2019
rect -31 -2053 -19 -2019
rect -77 -2059 -19 -2053
rect -77 -2127 -19 -2121
rect -77 -2161 -65 -2127
rect -31 -2161 -19 -2127
rect -77 -2167 -19 -2161
rect -119 -2220 -73 -2208
rect -119 -2796 -113 -2220
rect -79 -2796 -73 -2220
rect -119 -2808 -73 -2796
rect -23 -2220 23 -2208
rect -23 -2796 -17 -2220
rect 17 -2796 23 -2220
rect -23 -2808 23 -2796
rect 73 -2220 119 -2208
rect 73 -2796 79 -2220
rect 113 -2796 119 -2220
rect 73 -2808 119 -2796
rect 19 -2855 77 -2849
rect 19 -2889 31 -2855
rect 65 -2889 77 -2855
rect 19 -2895 77 -2889
rect 19 -2963 77 -2957
rect 19 -2997 31 -2963
rect 65 -2997 77 -2963
rect 19 -3003 77 -2997
rect -119 -3056 -73 -3044
rect -119 -3632 -113 -3056
rect -79 -3632 -73 -3056
rect -119 -3644 -73 -3632
rect -23 -3056 23 -3044
rect -23 -3632 -17 -3056
rect 17 -3632 23 -3056
rect -23 -3644 23 -3632
rect 73 -3056 119 -3044
rect 73 -3632 79 -3056
rect 113 -3632 119 -3056
rect 73 -3644 119 -3632
rect -77 -3691 -19 -3685
rect -77 -3725 -65 -3691
rect -31 -3725 -19 -3691
rect -77 -3731 -19 -3725
rect -77 -3799 -19 -3793
rect -77 -3833 -65 -3799
rect -31 -3833 -19 -3799
rect -77 -3839 -19 -3833
rect -119 -3892 -73 -3880
rect -119 -4468 -113 -3892
rect -79 -4468 -73 -3892
rect -119 -4480 -73 -4468
rect -23 -3892 23 -3880
rect -23 -4468 -17 -3892
rect 17 -4468 23 -3892
rect -23 -4480 23 -4468
rect 73 -3892 119 -3880
rect 73 -4468 79 -3892
rect 113 -4468 119 -3892
rect 73 -4480 119 -4468
rect 19 -4527 77 -4521
rect 19 -4561 31 -4527
rect 65 -4561 77 -4527
rect 19 -4567 77 -4561
rect 19 -4635 77 -4629
rect 19 -4669 31 -4635
rect 65 -4669 77 -4635
rect 19 -4675 77 -4669
rect -119 -4728 -73 -4716
rect -119 -5304 -113 -4728
rect -79 -5304 -73 -4728
rect -119 -5316 -73 -5304
rect -23 -4728 23 -4716
rect -23 -5304 -17 -4728
rect 17 -5304 23 -4728
rect -23 -5316 23 -5304
rect 73 -4728 119 -4716
rect 73 -5304 79 -4728
rect 113 -5304 119 -4728
rect 73 -5316 119 -5304
rect -77 -5363 -19 -5357
rect -77 -5397 -65 -5363
rect -31 -5397 -19 -5363
rect -77 -5403 -19 -5397
rect -77 -5471 -19 -5465
rect -77 -5505 -65 -5471
rect -31 -5505 -19 -5471
rect -77 -5511 -19 -5505
rect -119 -5564 -73 -5552
rect -119 -6140 -113 -5564
rect -79 -6140 -73 -5564
rect -119 -6152 -73 -6140
rect -23 -5564 23 -5552
rect -23 -6140 -17 -5564
rect 17 -6140 23 -5564
rect -23 -6152 23 -6140
rect 73 -5564 119 -5552
rect 73 -6140 79 -5564
rect 113 -6140 119 -5564
rect 73 -6152 119 -6140
rect 19 -6199 77 -6193
rect 19 -6233 31 -6199
rect 65 -6233 77 -6199
rect 19 -6239 77 -6233
rect 19 -6307 77 -6301
rect 19 -6341 31 -6307
rect 65 -6341 77 -6307
rect 19 -6347 77 -6341
rect -119 -6400 -73 -6388
rect -119 -6976 -113 -6400
rect -79 -6976 -73 -6400
rect -119 -6988 -73 -6976
rect -23 -6400 23 -6388
rect -23 -6976 -17 -6400
rect 17 -6976 23 -6400
rect -23 -6988 23 -6976
rect 73 -6400 119 -6388
rect 73 -6976 79 -6400
rect 113 -6976 119 -6400
rect 73 -6988 119 -6976
rect -77 -7035 -19 -7029
rect -77 -7069 -65 -7035
rect -31 -7069 -19 -7035
rect -77 -7075 -19 -7069
rect -77 -7143 -19 -7137
rect -77 -7177 -65 -7143
rect -31 -7177 -19 -7143
rect -77 -7183 -19 -7177
rect -119 -7236 -73 -7224
rect -119 -7812 -113 -7236
rect -79 -7812 -73 -7236
rect -119 -7824 -73 -7812
rect -23 -7236 23 -7224
rect -23 -7812 -17 -7236
rect 17 -7812 23 -7236
rect -23 -7824 23 -7812
rect 73 -7236 119 -7224
rect 73 -7812 79 -7236
rect 113 -7812 119 -7236
rect 73 -7824 119 -7812
rect 19 -7871 77 -7865
rect 19 -7905 31 -7871
rect 65 -7905 77 -7871
rect 19 -7911 77 -7905
rect 19 -7979 77 -7973
rect 19 -8013 31 -7979
rect 65 -8013 77 -7979
rect 19 -8019 77 -8013
rect -119 -8072 -73 -8060
rect -119 -8648 -113 -8072
rect -79 -8648 -73 -8072
rect -119 -8660 -73 -8648
rect -23 -8072 23 -8060
rect -23 -8648 -17 -8072
rect 17 -8648 23 -8072
rect -23 -8660 23 -8648
rect 73 -8072 119 -8060
rect 73 -8648 79 -8072
rect 113 -8648 119 -8072
rect 73 -8660 119 -8648
rect -77 -8707 -19 -8701
rect -77 -8741 -65 -8707
rect -31 -8741 -19 -8707
rect -77 -8747 -19 -8741
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -210 -8826 210 8826
string parameters w 3 l 0.15 m 21 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
