magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_p >>
rect -29 129 29 135
rect -29 95 -17 129
rect -29 89 29 95
<< nwell >>
rect -109 -182 109 148
<< pmos >>
rect -15 -120 15 48
<< pdiff >>
rect -73 15 -15 48
rect -73 -19 -61 15
rect -27 -19 -15 15
rect -73 -53 -15 -19
rect -73 -87 -61 -53
rect -27 -87 -15 -53
rect -73 -120 -15 -87
rect 15 15 73 48
rect 15 -19 27 15
rect 61 -19 73 15
rect 15 -53 73 -19
rect 15 -87 27 -53
rect 61 -87 73 -53
rect 15 -120 73 -87
<< pdiffc >>
rect -61 -19 -27 15
rect -61 -87 -27 -53
rect 27 -19 61 15
rect 27 -87 61 -53
<< poly >>
rect -33 129 33 145
rect -33 95 -17 129
rect 17 95 33 129
rect -33 79 33 95
rect -15 48 15 79
rect -15 -146 15 -120
<< polycont >>
rect -17 95 17 129
<< locali >>
rect -33 95 -17 129
rect 17 95 33 129
rect -61 17 -27 52
rect -61 -53 -27 -19
rect -61 -124 -27 -89
rect 27 17 61 52
rect 27 -53 61 -19
rect 27 -124 61 -89
<< viali >>
rect -17 95 17 129
rect -61 15 -27 17
rect -61 -17 -27 15
rect -61 -87 -27 -55
rect -61 -89 -27 -87
rect 27 15 61 17
rect 27 -17 61 15
rect 27 -87 61 -55
rect 27 -89 61 -87
<< metal1 >>
rect -29 129 29 135
rect -29 95 -17 129
rect 17 95 29 129
rect -29 89 29 95
rect -67 17 -21 48
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -55 -21 -17
rect -67 -89 -61 -55
rect -27 -89 -21 -55
rect -67 -120 -21 -89
rect 21 17 67 48
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -55 67 -17
rect 21 -89 27 -55
rect 61 -89 67 -55
rect 21 -120 67 -89
<< end >>
