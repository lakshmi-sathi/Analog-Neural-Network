magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< poly >>
rect 3963 675 4060 701
rect 3967 671 4060 675
rect 4030 623 4060 671
<< locali >>
rect 50 -150 4114 -118
rect 50 -184 85 -150
rect 119 -184 157 -150
rect 191 -184 229 -150
rect 263 -184 301 -150
rect 335 -184 373 -150
rect 407 -184 445 -150
rect 479 -184 517 -150
rect 551 -184 589 -150
rect 623 -184 661 -150
rect 695 -184 733 -150
rect 767 -184 805 -150
rect 839 -184 877 -150
rect 911 -184 949 -150
rect 983 -184 1021 -150
rect 1055 -184 1093 -150
rect 1127 -184 1165 -150
rect 1199 -184 1237 -150
rect 1271 -184 1309 -150
rect 1343 -184 1381 -150
rect 1415 -184 1453 -150
rect 1487 -184 1525 -150
rect 1559 -184 1597 -150
rect 1631 -184 1669 -150
rect 1703 -184 1741 -150
rect 1775 -184 1813 -150
rect 1847 -184 1885 -150
rect 1919 -184 1957 -150
rect 1991 -184 2029 -150
rect 2063 -184 2101 -150
rect 2135 -184 2173 -150
rect 2207 -184 2245 -150
rect 2279 -184 2317 -150
rect 2351 -184 2389 -150
rect 2423 -184 2461 -150
rect 2495 -184 2533 -150
rect 2567 -184 2605 -150
rect 2639 -184 2677 -150
rect 2711 -184 2749 -150
rect 2783 -184 2821 -150
rect 2855 -184 2893 -150
rect 2927 -184 2965 -150
rect 2999 -184 3037 -150
rect 3071 -184 3109 -150
rect 3143 -184 3181 -150
rect 3215 -184 3253 -150
rect 3287 -184 3325 -150
rect 3359 -184 3397 -150
rect 3431 -184 3469 -150
rect 3503 -184 3541 -150
rect 3575 -184 3613 -150
rect 3647 -184 3685 -150
rect 3719 -184 3757 -150
rect 3791 -184 3829 -150
rect 3863 -184 3901 -150
rect 3935 -184 3973 -150
rect 4007 -184 4045 -150
rect 4079 -184 4114 -150
rect 50 -216 4114 -184
<< viali >>
rect 85 -184 119 -150
rect 157 -184 191 -150
rect 229 -184 263 -150
rect 301 -184 335 -150
rect 373 -184 407 -150
rect 445 -184 479 -150
rect 517 -184 551 -150
rect 589 -184 623 -150
rect 661 -184 695 -150
rect 733 -184 767 -150
rect 805 -184 839 -150
rect 877 -184 911 -150
rect 949 -184 983 -150
rect 1021 -184 1055 -150
rect 1093 -184 1127 -150
rect 1165 -184 1199 -150
rect 1237 -184 1271 -150
rect 1309 -184 1343 -150
rect 1381 -184 1415 -150
rect 1453 -184 1487 -150
rect 1525 -184 1559 -150
rect 1597 -184 1631 -150
rect 1669 -184 1703 -150
rect 1741 -184 1775 -150
rect 1813 -184 1847 -150
rect 1885 -184 1919 -150
rect 1957 -184 1991 -150
rect 2029 -184 2063 -150
rect 2101 -184 2135 -150
rect 2173 -184 2207 -150
rect 2245 -184 2279 -150
rect 2317 -184 2351 -150
rect 2389 -184 2423 -150
rect 2461 -184 2495 -150
rect 2533 -184 2567 -150
rect 2605 -184 2639 -150
rect 2677 -184 2711 -150
rect 2749 -184 2783 -150
rect 2821 -184 2855 -150
rect 2893 -184 2927 -150
rect 2965 -184 2999 -150
rect 3037 -184 3071 -150
rect 3109 -184 3143 -150
rect 3181 -184 3215 -150
rect 3253 -184 3287 -150
rect 3325 -184 3359 -150
rect 3397 -184 3431 -150
rect 3469 -184 3503 -150
rect 3541 -184 3575 -150
rect 3613 -184 3647 -150
rect 3685 -184 3719 -150
rect 3757 -184 3791 -150
rect 3829 -184 3863 -150
rect 3901 -184 3935 -150
rect 3973 -184 4007 -150
rect 4045 -184 4079 -150
<< metal1 >>
rect 76 654 3980 706
rect 126 620 188 622
rect 318 620 380 622
rect 510 620 572 622
rect 702 620 764 622
rect 894 620 956 622
rect 1086 620 1148 622
rect 1278 620 1340 622
rect 1470 620 1532 622
rect 1662 620 1724 622
rect 1854 620 1916 622
rect 2046 620 2108 622
rect 2238 620 2300 622
rect 2430 620 2492 622
rect 2622 620 2684 622
rect 2814 620 2876 622
rect 3006 620 3068 622
rect 3198 620 3260 622
rect 3390 620 3452 622
rect 3582 620 3644 622
rect 3774 620 3836 622
rect 3966 620 4028 622
rect 126 611 190 620
rect 126 559 132 611
rect 184 559 190 611
rect 126 547 190 559
rect 126 495 132 547
rect 184 495 190 547
rect 126 483 190 495
rect 126 431 132 483
rect 184 431 190 483
rect 126 419 190 431
rect 126 367 132 419
rect 184 367 190 419
rect 126 364 190 367
rect 318 611 382 620
rect 318 559 324 611
rect 376 559 382 611
rect 318 547 382 559
rect 318 495 324 547
rect 376 495 382 547
rect 318 483 382 495
rect 318 431 324 483
rect 376 431 382 483
rect 318 419 382 431
rect 318 367 324 419
rect 376 367 382 419
rect 318 364 382 367
rect 510 611 574 620
rect 510 559 516 611
rect 568 559 574 611
rect 510 547 574 559
rect 510 495 516 547
rect 568 495 574 547
rect 510 483 574 495
rect 510 431 516 483
rect 568 431 574 483
rect 510 419 574 431
rect 510 367 516 419
rect 568 367 574 419
rect 510 364 574 367
rect 702 611 766 620
rect 702 559 708 611
rect 760 559 766 611
rect 702 547 766 559
rect 702 495 708 547
rect 760 495 766 547
rect 702 483 766 495
rect 702 431 708 483
rect 760 431 766 483
rect 702 419 766 431
rect 702 367 708 419
rect 760 367 766 419
rect 702 364 766 367
rect 894 611 958 620
rect 894 559 900 611
rect 952 559 958 611
rect 894 547 958 559
rect 894 495 900 547
rect 952 495 958 547
rect 894 483 958 495
rect 894 431 900 483
rect 952 431 958 483
rect 894 419 958 431
rect 894 367 900 419
rect 952 367 958 419
rect 894 364 958 367
rect 1086 611 1150 620
rect 1086 559 1092 611
rect 1144 559 1150 611
rect 1086 547 1150 559
rect 1086 495 1092 547
rect 1144 495 1150 547
rect 1086 483 1150 495
rect 1086 431 1092 483
rect 1144 431 1150 483
rect 1086 419 1150 431
rect 1086 367 1092 419
rect 1144 367 1150 419
rect 1086 364 1150 367
rect 1278 611 1342 620
rect 1278 559 1284 611
rect 1336 559 1342 611
rect 1278 547 1342 559
rect 1278 495 1284 547
rect 1336 495 1342 547
rect 1278 483 1342 495
rect 1278 431 1284 483
rect 1336 431 1342 483
rect 1278 419 1342 431
rect 1278 367 1284 419
rect 1336 367 1342 419
rect 1278 364 1342 367
rect 1470 611 1534 620
rect 1470 559 1476 611
rect 1528 559 1534 611
rect 1470 547 1534 559
rect 1470 495 1476 547
rect 1528 495 1534 547
rect 1470 483 1534 495
rect 1470 431 1476 483
rect 1528 431 1534 483
rect 1470 419 1534 431
rect 1470 367 1476 419
rect 1528 367 1534 419
rect 1470 364 1534 367
rect 1662 611 1726 620
rect 1662 559 1668 611
rect 1720 559 1726 611
rect 1662 547 1726 559
rect 1662 495 1668 547
rect 1720 495 1726 547
rect 1662 483 1726 495
rect 1662 431 1668 483
rect 1720 431 1726 483
rect 1662 419 1726 431
rect 1662 367 1668 419
rect 1720 367 1726 419
rect 1662 364 1726 367
rect 1854 611 1918 620
rect 1854 559 1860 611
rect 1912 559 1918 611
rect 1854 547 1918 559
rect 1854 495 1860 547
rect 1912 495 1918 547
rect 1854 483 1918 495
rect 1854 431 1860 483
rect 1912 431 1918 483
rect 1854 419 1918 431
rect 1854 367 1860 419
rect 1912 367 1918 419
rect 1854 364 1918 367
rect 2046 611 2110 620
rect 2046 559 2052 611
rect 2104 559 2110 611
rect 2046 547 2110 559
rect 2046 495 2052 547
rect 2104 495 2110 547
rect 2046 483 2110 495
rect 2046 431 2052 483
rect 2104 431 2110 483
rect 2046 419 2110 431
rect 2046 367 2052 419
rect 2104 367 2110 419
rect 2046 364 2110 367
rect 2238 611 2302 620
rect 2238 559 2244 611
rect 2296 559 2302 611
rect 2238 547 2302 559
rect 2238 495 2244 547
rect 2296 495 2302 547
rect 2238 483 2302 495
rect 2238 431 2244 483
rect 2296 431 2302 483
rect 2238 419 2302 431
rect 2238 367 2244 419
rect 2296 367 2302 419
rect 2238 364 2302 367
rect 2430 611 2494 620
rect 2430 559 2436 611
rect 2488 559 2494 611
rect 2430 547 2494 559
rect 2430 495 2436 547
rect 2488 495 2494 547
rect 2430 483 2494 495
rect 2430 431 2436 483
rect 2488 431 2494 483
rect 2430 419 2494 431
rect 2430 367 2436 419
rect 2488 367 2494 419
rect 2430 364 2494 367
rect 2622 611 2686 620
rect 2622 559 2628 611
rect 2680 559 2686 611
rect 2622 547 2686 559
rect 2622 495 2628 547
rect 2680 495 2686 547
rect 2622 483 2686 495
rect 2622 431 2628 483
rect 2680 431 2686 483
rect 2622 419 2686 431
rect 2622 367 2628 419
rect 2680 367 2686 419
rect 2622 364 2686 367
rect 2814 611 2878 620
rect 2814 559 2820 611
rect 2872 559 2878 611
rect 2814 547 2878 559
rect 2814 495 2820 547
rect 2872 495 2878 547
rect 2814 483 2878 495
rect 2814 431 2820 483
rect 2872 431 2878 483
rect 2814 419 2878 431
rect 2814 367 2820 419
rect 2872 367 2878 419
rect 2814 364 2878 367
rect 3006 611 3070 620
rect 3006 559 3012 611
rect 3064 559 3070 611
rect 3006 547 3070 559
rect 3006 495 3012 547
rect 3064 495 3070 547
rect 3006 483 3070 495
rect 3006 431 3012 483
rect 3064 431 3070 483
rect 3006 419 3070 431
rect 3006 367 3012 419
rect 3064 367 3070 419
rect 3006 364 3070 367
rect 3198 611 3262 620
rect 3198 559 3204 611
rect 3256 559 3262 611
rect 3198 547 3262 559
rect 3198 495 3204 547
rect 3256 495 3262 547
rect 3198 483 3262 495
rect 3198 431 3204 483
rect 3256 431 3262 483
rect 3198 419 3262 431
rect 3198 367 3204 419
rect 3256 367 3262 419
rect 3198 364 3262 367
rect 3390 611 3454 620
rect 3390 559 3396 611
rect 3448 559 3454 611
rect 3390 547 3454 559
rect 3390 495 3396 547
rect 3448 495 3454 547
rect 3390 483 3454 495
rect 3390 431 3396 483
rect 3448 431 3454 483
rect 3390 419 3454 431
rect 3390 367 3396 419
rect 3448 367 3454 419
rect 3390 364 3454 367
rect 3582 611 3646 620
rect 3582 559 3588 611
rect 3640 559 3646 611
rect 3582 547 3646 559
rect 3582 495 3588 547
rect 3640 495 3646 547
rect 3582 483 3646 495
rect 3582 431 3588 483
rect 3640 431 3646 483
rect 3582 419 3646 431
rect 3582 367 3588 419
rect 3640 367 3646 419
rect 3582 364 3646 367
rect 3774 611 3838 620
rect 3774 559 3780 611
rect 3832 559 3838 611
rect 3774 547 3838 559
rect 3774 495 3780 547
rect 3832 495 3838 547
rect 3774 483 3838 495
rect 3774 431 3780 483
rect 3832 431 3838 483
rect 3774 419 3838 431
rect 3774 367 3780 419
rect 3832 367 3838 419
rect 3774 364 3838 367
rect 3966 611 4030 620
rect 3966 559 3972 611
rect 4024 559 4030 611
rect 3966 547 4030 559
rect 3966 495 3972 547
rect 4024 495 4030 547
rect 3966 483 4030 495
rect 3966 431 3972 483
rect 4024 431 4030 483
rect 3966 419 4030 431
rect 3966 367 3972 419
rect 4024 367 4030 419
rect 3966 364 4030 367
rect 30 279 94 284
rect 30 227 36 279
rect 88 227 94 279
rect 30 215 94 227
rect 30 163 36 215
rect 88 163 94 215
rect 30 151 94 163
rect 30 99 36 151
rect 88 99 94 151
rect 30 87 94 99
rect 30 35 36 87
rect 88 35 94 87
rect 30 24 94 35
rect 222 279 286 284
rect 222 227 228 279
rect 280 227 286 279
rect 222 215 286 227
rect 222 163 228 215
rect 280 163 286 215
rect 222 151 286 163
rect 222 99 228 151
rect 280 99 286 151
rect 222 87 286 99
rect 222 35 228 87
rect 280 35 286 87
rect 222 24 286 35
rect 414 279 478 284
rect 414 227 420 279
rect 472 227 478 279
rect 414 215 478 227
rect 414 163 420 215
rect 472 163 478 215
rect 414 151 478 163
rect 414 99 420 151
rect 472 99 478 151
rect 414 87 478 99
rect 414 35 420 87
rect 472 35 478 87
rect 414 24 478 35
rect 606 279 670 284
rect 606 227 612 279
rect 664 227 670 279
rect 606 215 670 227
rect 606 163 612 215
rect 664 163 670 215
rect 606 151 670 163
rect 606 99 612 151
rect 664 99 670 151
rect 606 87 670 99
rect 606 35 612 87
rect 664 35 670 87
rect 606 24 670 35
rect 798 279 862 284
rect 798 227 804 279
rect 856 227 862 279
rect 798 215 862 227
rect 798 163 804 215
rect 856 163 862 215
rect 798 151 862 163
rect 798 99 804 151
rect 856 99 862 151
rect 798 87 862 99
rect 798 35 804 87
rect 856 35 862 87
rect 798 24 862 35
rect 990 279 1054 284
rect 990 227 996 279
rect 1048 227 1054 279
rect 990 215 1054 227
rect 990 163 996 215
rect 1048 163 1054 215
rect 990 151 1054 163
rect 990 99 996 151
rect 1048 99 1054 151
rect 990 87 1054 99
rect 990 35 996 87
rect 1048 35 1054 87
rect 990 24 1054 35
rect 1182 279 1246 284
rect 1182 227 1188 279
rect 1240 227 1246 279
rect 1182 215 1246 227
rect 1182 163 1188 215
rect 1240 163 1246 215
rect 1182 151 1246 163
rect 1182 99 1188 151
rect 1240 99 1246 151
rect 1182 87 1246 99
rect 1182 35 1188 87
rect 1240 35 1246 87
rect 1182 24 1246 35
rect 1374 279 1438 284
rect 1374 227 1380 279
rect 1432 227 1438 279
rect 1374 215 1438 227
rect 1374 163 1380 215
rect 1432 163 1438 215
rect 1374 151 1438 163
rect 1374 99 1380 151
rect 1432 99 1438 151
rect 1374 87 1438 99
rect 1374 35 1380 87
rect 1432 35 1438 87
rect 1374 24 1438 35
rect 1566 279 1630 284
rect 1566 227 1572 279
rect 1624 227 1630 279
rect 1566 215 1630 227
rect 1566 163 1572 215
rect 1624 163 1630 215
rect 1566 151 1630 163
rect 1566 99 1572 151
rect 1624 99 1630 151
rect 1566 87 1630 99
rect 1566 35 1572 87
rect 1624 35 1630 87
rect 1566 24 1630 35
rect 1758 279 1822 284
rect 1758 227 1764 279
rect 1816 227 1822 279
rect 1758 215 1822 227
rect 1758 163 1764 215
rect 1816 163 1822 215
rect 1758 151 1822 163
rect 1758 99 1764 151
rect 1816 99 1822 151
rect 1758 87 1822 99
rect 1758 35 1764 87
rect 1816 35 1822 87
rect 1758 24 1822 35
rect 1950 279 2014 284
rect 1950 227 1956 279
rect 2008 227 2014 279
rect 1950 215 2014 227
rect 1950 163 1956 215
rect 2008 163 2014 215
rect 1950 151 2014 163
rect 1950 99 1956 151
rect 2008 99 2014 151
rect 1950 87 2014 99
rect 1950 35 1956 87
rect 2008 35 2014 87
rect 1950 24 2014 35
rect 2142 279 2206 284
rect 2142 227 2148 279
rect 2200 227 2206 279
rect 2142 215 2206 227
rect 2142 163 2148 215
rect 2200 163 2206 215
rect 2142 151 2206 163
rect 2142 99 2148 151
rect 2200 99 2206 151
rect 2142 87 2206 99
rect 2142 35 2148 87
rect 2200 35 2206 87
rect 2142 24 2206 35
rect 2334 279 2398 284
rect 2334 227 2340 279
rect 2392 227 2398 279
rect 2334 215 2398 227
rect 2334 163 2340 215
rect 2392 163 2398 215
rect 2334 151 2398 163
rect 2334 99 2340 151
rect 2392 99 2398 151
rect 2334 87 2398 99
rect 2334 35 2340 87
rect 2392 35 2398 87
rect 2334 24 2398 35
rect 2526 279 2590 284
rect 2526 227 2532 279
rect 2584 227 2590 279
rect 2526 215 2590 227
rect 2526 163 2532 215
rect 2584 163 2590 215
rect 2526 151 2590 163
rect 2526 99 2532 151
rect 2584 99 2590 151
rect 2526 87 2590 99
rect 2526 35 2532 87
rect 2584 35 2590 87
rect 2526 24 2590 35
rect 2718 279 2782 284
rect 2718 227 2724 279
rect 2776 227 2782 279
rect 2718 215 2782 227
rect 2718 163 2724 215
rect 2776 163 2782 215
rect 2718 151 2782 163
rect 2718 99 2724 151
rect 2776 99 2782 151
rect 2718 87 2782 99
rect 2718 35 2724 87
rect 2776 35 2782 87
rect 2718 24 2782 35
rect 2910 279 2974 284
rect 2910 227 2916 279
rect 2968 227 2974 279
rect 2910 215 2974 227
rect 2910 163 2916 215
rect 2968 163 2974 215
rect 2910 151 2974 163
rect 2910 99 2916 151
rect 2968 99 2974 151
rect 2910 87 2974 99
rect 2910 35 2916 87
rect 2968 35 2974 87
rect 2910 24 2974 35
rect 3102 279 3166 284
rect 3102 227 3108 279
rect 3160 227 3166 279
rect 3102 215 3166 227
rect 3102 163 3108 215
rect 3160 163 3166 215
rect 3102 151 3166 163
rect 3102 99 3108 151
rect 3160 99 3166 151
rect 3102 87 3166 99
rect 3102 35 3108 87
rect 3160 35 3166 87
rect 3102 24 3166 35
rect 3294 279 3358 284
rect 3294 227 3300 279
rect 3352 227 3358 279
rect 3294 215 3358 227
rect 3294 163 3300 215
rect 3352 163 3358 215
rect 3294 151 3358 163
rect 3294 99 3300 151
rect 3352 99 3358 151
rect 3294 87 3358 99
rect 3294 35 3300 87
rect 3352 35 3358 87
rect 3294 24 3358 35
rect 3486 279 3550 284
rect 3486 227 3492 279
rect 3544 227 3550 279
rect 3486 215 3550 227
rect 3486 163 3492 215
rect 3544 163 3550 215
rect 3486 151 3550 163
rect 3486 99 3492 151
rect 3544 99 3550 151
rect 3486 87 3550 99
rect 3486 35 3492 87
rect 3544 35 3550 87
rect 3486 24 3550 35
rect 3678 279 3742 284
rect 3678 227 3684 279
rect 3736 227 3742 279
rect 3678 215 3742 227
rect 3678 163 3684 215
rect 3736 163 3742 215
rect 3678 151 3742 163
rect 3678 99 3684 151
rect 3736 99 3742 151
rect 3678 87 3742 99
rect 3678 35 3684 87
rect 3736 35 3742 87
rect 3678 24 3742 35
rect 3870 279 3934 284
rect 3870 227 3876 279
rect 3928 227 3934 279
rect 3870 215 3934 227
rect 3870 163 3876 215
rect 3928 163 3934 215
rect 3870 151 3934 163
rect 3870 99 3876 151
rect 3928 99 3934 151
rect 3870 87 3934 99
rect 3870 35 3876 87
rect 3928 35 3934 87
rect 3870 24 3934 35
rect 4062 279 4126 284
rect 4062 227 4068 279
rect 4120 227 4126 279
rect 4062 215 4126 227
rect 4062 163 4068 215
rect 4120 163 4126 215
rect 4062 151 4126 163
rect 4062 99 4068 151
rect 4120 99 4126 151
rect 4062 87 4126 99
rect 4062 35 4068 87
rect 4120 35 4126 87
rect 4062 24 4126 35
rect 172 -60 4076 -8
rect 50 -142 4114 -116
rect 50 -194 73 -142
rect 125 -194 137 -142
rect 189 -150 201 -142
rect 253 -150 265 -142
rect 317 -150 329 -142
rect 381 -150 393 -142
rect 445 -150 457 -142
rect 509 -150 521 -142
rect 191 -184 201 -150
rect 263 -184 265 -150
rect 509 -184 517 -150
rect 189 -194 201 -184
rect 253 -194 265 -184
rect 317 -194 329 -184
rect 381 -194 393 -184
rect 445 -194 457 -184
rect 509 -194 521 -184
rect 573 -194 585 -142
rect 637 -194 649 -142
rect 701 -194 713 -142
rect 765 -150 777 -142
rect 829 -150 841 -142
rect 893 -150 905 -142
rect 957 -150 969 -142
rect 1021 -150 1033 -142
rect 1085 -150 1097 -142
rect 767 -184 777 -150
rect 839 -184 841 -150
rect 1085 -184 1093 -150
rect 765 -194 777 -184
rect 829 -194 841 -184
rect 893 -194 905 -184
rect 957 -194 969 -184
rect 1021 -194 1033 -184
rect 1085 -194 1097 -184
rect 1149 -194 1161 -142
rect 1213 -194 1225 -142
rect 1277 -194 1289 -142
rect 1341 -150 1353 -142
rect 1405 -150 1417 -142
rect 1469 -150 1481 -142
rect 1533 -150 1545 -142
rect 1597 -150 1609 -142
rect 1661 -150 1673 -142
rect 1343 -184 1353 -150
rect 1415 -184 1417 -150
rect 1661 -184 1669 -150
rect 1341 -194 1353 -184
rect 1405 -194 1417 -184
rect 1469 -194 1481 -184
rect 1533 -194 1545 -184
rect 1597 -194 1609 -184
rect 1661 -194 1673 -184
rect 1725 -194 1737 -142
rect 1789 -194 1801 -142
rect 1853 -194 1865 -142
rect 1917 -150 1929 -142
rect 1981 -150 1993 -142
rect 2045 -150 2057 -142
rect 2109 -150 2121 -142
rect 2173 -150 2185 -142
rect 2237 -150 2249 -142
rect 1919 -184 1929 -150
rect 1991 -184 1993 -150
rect 2237 -184 2245 -150
rect 1917 -194 1929 -184
rect 1981 -194 1993 -184
rect 2045 -194 2057 -184
rect 2109 -194 2121 -184
rect 2173 -194 2185 -184
rect 2237 -194 2249 -184
rect 2301 -194 2313 -142
rect 2365 -194 2377 -142
rect 2429 -194 2441 -142
rect 2493 -150 2505 -142
rect 2557 -150 2569 -142
rect 2621 -150 2633 -142
rect 2685 -150 2697 -142
rect 2749 -150 2761 -142
rect 2813 -150 2825 -142
rect 2495 -184 2505 -150
rect 2567 -184 2569 -150
rect 2813 -184 2821 -150
rect 2493 -194 2505 -184
rect 2557 -194 2569 -184
rect 2621 -194 2633 -184
rect 2685 -194 2697 -184
rect 2749 -194 2761 -184
rect 2813 -194 2825 -184
rect 2877 -194 2889 -142
rect 2941 -194 2953 -142
rect 3005 -194 3017 -142
rect 3069 -150 3081 -142
rect 3133 -150 3145 -142
rect 3197 -150 3209 -142
rect 3261 -150 3273 -142
rect 3325 -150 3337 -142
rect 3389 -150 3401 -142
rect 3071 -184 3081 -150
rect 3143 -184 3145 -150
rect 3389 -184 3397 -150
rect 3069 -194 3081 -184
rect 3133 -194 3145 -184
rect 3197 -194 3209 -184
rect 3261 -194 3273 -184
rect 3325 -194 3337 -184
rect 3389 -194 3401 -184
rect 3453 -194 3465 -142
rect 3517 -194 3529 -142
rect 3581 -194 3593 -142
rect 3645 -150 3657 -142
rect 3709 -150 3721 -142
rect 3773 -150 3785 -142
rect 3837 -150 3849 -142
rect 3901 -150 3913 -142
rect 3965 -150 3977 -142
rect 3647 -184 3657 -150
rect 3719 -184 3721 -150
rect 3965 -184 3973 -150
rect 3645 -194 3657 -184
rect 3709 -194 3721 -184
rect 3773 -194 3785 -184
rect 3837 -194 3849 -184
rect 3901 -194 3913 -184
rect 3965 -194 3977 -184
rect 4029 -194 4041 -142
rect 4093 -194 4114 -142
rect 50 -220 4114 -194
<< via1 >>
rect 132 559 184 611
rect 132 495 184 547
rect 132 431 184 483
rect 132 367 184 419
rect 324 559 376 611
rect 324 495 376 547
rect 324 431 376 483
rect 324 367 376 419
rect 516 559 568 611
rect 516 495 568 547
rect 516 431 568 483
rect 516 367 568 419
rect 708 559 760 611
rect 708 495 760 547
rect 708 431 760 483
rect 708 367 760 419
rect 900 559 952 611
rect 900 495 952 547
rect 900 431 952 483
rect 900 367 952 419
rect 1092 559 1144 611
rect 1092 495 1144 547
rect 1092 431 1144 483
rect 1092 367 1144 419
rect 1284 559 1336 611
rect 1284 495 1336 547
rect 1284 431 1336 483
rect 1284 367 1336 419
rect 1476 559 1528 611
rect 1476 495 1528 547
rect 1476 431 1528 483
rect 1476 367 1528 419
rect 1668 559 1720 611
rect 1668 495 1720 547
rect 1668 431 1720 483
rect 1668 367 1720 419
rect 1860 559 1912 611
rect 1860 495 1912 547
rect 1860 431 1912 483
rect 1860 367 1912 419
rect 2052 559 2104 611
rect 2052 495 2104 547
rect 2052 431 2104 483
rect 2052 367 2104 419
rect 2244 559 2296 611
rect 2244 495 2296 547
rect 2244 431 2296 483
rect 2244 367 2296 419
rect 2436 559 2488 611
rect 2436 495 2488 547
rect 2436 431 2488 483
rect 2436 367 2488 419
rect 2628 559 2680 611
rect 2628 495 2680 547
rect 2628 431 2680 483
rect 2628 367 2680 419
rect 2820 559 2872 611
rect 2820 495 2872 547
rect 2820 431 2872 483
rect 2820 367 2872 419
rect 3012 559 3064 611
rect 3012 495 3064 547
rect 3012 431 3064 483
rect 3012 367 3064 419
rect 3204 559 3256 611
rect 3204 495 3256 547
rect 3204 431 3256 483
rect 3204 367 3256 419
rect 3396 559 3448 611
rect 3396 495 3448 547
rect 3396 431 3448 483
rect 3396 367 3448 419
rect 3588 559 3640 611
rect 3588 495 3640 547
rect 3588 431 3640 483
rect 3588 367 3640 419
rect 3780 559 3832 611
rect 3780 495 3832 547
rect 3780 431 3832 483
rect 3780 367 3832 419
rect 3972 559 4024 611
rect 3972 495 4024 547
rect 3972 431 4024 483
rect 3972 367 4024 419
rect 36 227 88 279
rect 36 163 88 215
rect 36 99 88 151
rect 36 35 88 87
rect 228 227 280 279
rect 228 163 280 215
rect 228 99 280 151
rect 228 35 280 87
rect 420 227 472 279
rect 420 163 472 215
rect 420 99 472 151
rect 420 35 472 87
rect 612 227 664 279
rect 612 163 664 215
rect 612 99 664 151
rect 612 35 664 87
rect 804 227 856 279
rect 804 163 856 215
rect 804 99 856 151
rect 804 35 856 87
rect 996 227 1048 279
rect 996 163 1048 215
rect 996 99 1048 151
rect 996 35 1048 87
rect 1188 227 1240 279
rect 1188 163 1240 215
rect 1188 99 1240 151
rect 1188 35 1240 87
rect 1380 227 1432 279
rect 1380 163 1432 215
rect 1380 99 1432 151
rect 1380 35 1432 87
rect 1572 227 1624 279
rect 1572 163 1624 215
rect 1572 99 1624 151
rect 1572 35 1624 87
rect 1764 227 1816 279
rect 1764 163 1816 215
rect 1764 99 1816 151
rect 1764 35 1816 87
rect 1956 227 2008 279
rect 1956 163 2008 215
rect 1956 99 2008 151
rect 1956 35 2008 87
rect 2148 227 2200 279
rect 2148 163 2200 215
rect 2148 99 2200 151
rect 2148 35 2200 87
rect 2340 227 2392 279
rect 2340 163 2392 215
rect 2340 99 2392 151
rect 2340 35 2392 87
rect 2532 227 2584 279
rect 2532 163 2584 215
rect 2532 99 2584 151
rect 2532 35 2584 87
rect 2724 227 2776 279
rect 2724 163 2776 215
rect 2724 99 2776 151
rect 2724 35 2776 87
rect 2916 227 2968 279
rect 2916 163 2968 215
rect 2916 99 2968 151
rect 2916 35 2968 87
rect 3108 227 3160 279
rect 3108 163 3160 215
rect 3108 99 3160 151
rect 3108 35 3160 87
rect 3300 227 3352 279
rect 3300 163 3352 215
rect 3300 99 3352 151
rect 3300 35 3352 87
rect 3492 227 3544 279
rect 3492 163 3544 215
rect 3492 99 3544 151
rect 3492 35 3544 87
rect 3684 227 3736 279
rect 3684 163 3736 215
rect 3684 99 3736 151
rect 3684 35 3736 87
rect 3876 227 3928 279
rect 3876 163 3928 215
rect 3876 99 3928 151
rect 3876 35 3928 87
rect 4068 227 4120 279
rect 4068 163 4120 215
rect 4068 99 4120 151
rect 4068 35 4120 87
rect 73 -150 125 -142
rect 73 -184 85 -150
rect 85 -184 119 -150
rect 119 -184 125 -150
rect 73 -194 125 -184
rect 137 -150 189 -142
rect 201 -150 253 -142
rect 265 -150 317 -142
rect 329 -150 381 -142
rect 393 -150 445 -142
rect 457 -150 509 -142
rect 521 -150 573 -142
rect 137 -184 157 -150
rect 157 -184 189 -150
rect 201 -184 229 -150
rect 229 -184 253 -150
rect 265 -184 301 -150
rect 301 -184 317 -150
rect 329 -184 335 -150
rect 335 -184 373 -150
rect 373 -184 381 -150
rect 393 -184 407 -150
rect 407 -184 445 -150
rect 457 -184 479 -150
rect 479 -184 509 -150
rect 521 -184 551 -150
rect 551 -184 573 -150
rect 137 -194 189 -184
rect 201 -194 253 -184
rect 265 -194 317 -184
rect 329 -194 381 -184
rect 393 -194 445 -184
rect 457 -194 509 -184
rect 521 -194 573 -184
rect 585 -150 637 -142
rect 585 -184 589 -150
rect 589 -184 623 -150
rect 623 -184 637 -150
rect 585 -194 637 -184
rect 649 -150 701 -142
rect 649 -184 661 -150
rect 661 -184 695 -150
rect 695 -184 701 -150
rect 649 -194 701 -184
rect 713 -150 765 -142
rect 777 -150 829 -142
rect 841 -150 893 -142
rect 905 -150 957 -142
rect 969 -150 1021 -142
rect 1033 -150 1085 -142
rect 1097 -150 1149 -142
rect 713 -184 733 -150
rect 733 -184 765 -150
rect 777 -184 805 -150
rect 805 -184 829 -150
rect 841 -184 877 -150
rect 877 -184 893 -150
rect 905 -184 911 -150
rect 911 -184 949 -150
rect 949 -184 957 -150
rect 969 -184 983 -150
rect 983 -184 1021 -150
rect 1033 -184 1055 -150
rect 1055 -184 1085 -150
rect 1097 -184 1127 -150
rect 1127 -184 1149 -150
rect 713 -194 765 -184
rect 777 -194 829 -184
rect 841 -194 893 -184
rect 905 -194 957 -184
rect 969 -194 1021 -184
rect 1033 -194 1085 -184
rect 1097 -194 1149 -184
rect 1161 -150 1213 -142
rect 1161 -184 1165 -150
rect 1165 -184 1199 -150
rect 1199 -184 1213 -150
rect 1161 -194 1213 -184
rect 1225 -150 1277 -142
rect 1225 -184 1237 -150
rect 1237 -184 1271 -150
rect 1271 -184 1277 -150
rect 1225 -194 1277 -184
rect 1289 -150 1341 -142
rect 1353 -150 1405 -142
rect 1417 -150 1469 -142
rect 1481 -150 1533 -142
rect 1545 -150 1597 -142
rect 1609 -150 1661 -142
rect 1673 -150 1725 -142
rect 1289 -184 1309 -150
rect 1309 -184 1341 -150
rect 1353 -184 1381 -150
rect 1381 -184 1405 -150
rect 1417 -184 1453 -150
rect 1453 -184 1469 -150
rect 1481 -184 1487 -150
rect 1487 -184 1525 -150
rect 1525 -184 1533 -150
rect 1545 -184 1559 -150
rect 1559 -184 1597 -150
rect 1609 -184 1631 -150
rect 1631 -184 1661 -150
rect 1673 -184 1703 -150
rect 1703 -184 1725 -150
rect 1289 -194 1341 -184
rect 1353 -194 1405 -184
rect 1417 -194 1469 -184
rect 1481 -194 1533 -184
rect 1545 -194 1597 -184
rect 1609 -194 1661 -184
rect 1673 -194 1725 -184
rect 1737 -150 1789 -142
rect 1737 -184 1741 -150
rect 1741 -184 1775 -150
rect 1775 -184 1789 -150
rect 1737 -194 1789 -184
rect 1801 -150 1853 -142
rect 1801 -184 1813 -150
rect 1813 -184 1847 -150
rect 1847 -184 1853 -150
rect 1801 -194 1853 -184
rect 1865 -150 1917 -142
rect 1929 -150 1981 -142
rect 1993 -150 2045 -142
rect 2057 -150 2109 -142
rect 2121 -150 2173 -142
rect 2185 -150 2237 -142
rect 2249 -150 2301 -142
rect 1865 -184 1885 -150
rect 1885 -184 1917 -150
rect 1929 -184 1957 -150
rect 1957 -184 1981 -150
rect 1993 -184 2029 -150
rect 2029 -184 2045 -150
rect 2057 -184 2063 -150
rect 2063 -184 2101 -150
rect 2101 -184 2109 -150
rect 2121 -184 2135 -150
rect 2135 -184 2173 -150
rect 2185 -184 2207 -150
rect 2207 -184 2237 -150
rect 2249 -184 2279 -150
rect 2279 -184 2301 -150
rect 1865 -194 1917 -184
rect 1929 -194 1981 -184
rect 1993 -194 2045 -184
rect 2057 -194 2109 -184
rect 2121 -194 2173 -184
rect 2185 -194 2237 -184
rect 2249 -194 2301 -184
rect 2313 -150 2365 -142
rect 2313 -184 2317 -150
rect 2317 -184 2351 -150
rect 2351 -184 2365 -150
rect 2313 -194 2365 -184
rect 2377 -150 2429 -142
rect 2377 -184 2389 -150
rect 2389 -184 2423 -150
rect 2423 -184 2429 -150
rect 2377 -194 2429 -184
rect 2441 -150 2493 -142
rect 2505 -150 2557 -142
rect 2569 -150 2621 -142
rect 2633 -150 2685 -142
rect 2697 -150 2749 -142
rect 2761 -150 2813 -142
rect 2825 -150 2877 -142
rect 2441 -184 2461 -150
rect 2461 -184 2493 -150
rect 2505 -184 2533 -150
rect 2533 -184 2557 -150
rect 2569 -184 2605 -150
rect 2605 -184 2621 -150
rect 2633 -184 2639 -150
rect 2639 -184 2677 -150
rect 2677 -184 2685 -150
rect 2697 -184 2711 -150
rect 2711 -184 2749 -150
rect 2761 -184 2783 -150
rect 2783 -184 2813 -150
rect 2825 -184 2855 -150
rect 2855 -184 2877 -150
rect 2441 -194 2493 -184
rect 2505 -194 2557 -184
rect 2569 -194 2621 -184
rect 2633 -194 2685 -184
rect 2697 -194 2749 -184
rect 2761 -194 2813 -184
rect 2825 -194 2877 -184
rect 2889 -150 2941 -142
rect 2889 -184 2893 -150
rect 2893 -184 2927 -150
rect 2927 -184 2941 -150
rect 2889 -194 2941 -184
rect 2953 -150 3005 -142
rect 2953 -184 2965 -150
rect 2965 -184 2999 -150
rect 2999 -184 3005 -150
rect 2953 -194 3005 -184
rect 3017 -150 3069 -142
rect 3081 -150 3133 -142
rect 3145 -150 3197 -142
rect 3209 -150 3261 -142
rect 3273 -150 3325 -142
rect 3337 -150 3389 -142
rect 3401 -150 3453 -142
rect 3017 -184 3037 -150
rect 3037 -184 3069 -150
rect 3081 -184 3109 -150
rect 3109 -184 3133 -150
rect 3145 -184 3181 -150
rect 3181 -184 3197 -150
rect 3209 -184 3215 -150
rect 3215 -184 3253 -150
rect 3253 -184 3261 -150
rect 3273 -184 3287 -150
rect 3287 -184 3325 -150
rect 3337 -184 3359 -150
rect 3359 -184 3389 -150
rect 3401 -184 3431 -150
rect 3431 -184 3453 -150
rect 3017 -194 3069 -184
rect 3081 -194 3133 -184
rect 3145 -194 3197 -184
rect 3209 -194 3261 -184
rect 3273 -194 3325 -184
rect 3337 -194 3389 -184
rect 3401 -194 3453 -184
rect 3465 -150 3517 -142
rect 3465 -184 3469 -150
rect 3469 -184 3503 -150
rect 3503 -184 3517 -150
rect 3465 -194 3517 -184
rect 3529 -150 3581 -142
rect 3529 -184 3541 -150
rect 3541 -184 3575 -150
rect 3575 -184 3581 -150
rect 3529 -194 3581 -184
rect 3593 -150 3645 -142
rect 3657 -150 3709 -142
rect 3721 -150 3773 -142
rect 3785 -150 3837 -142
rect 3849 -150 3901 -142
rect 3913 -150 3965 -142
rect 3977 -150 4029 -142
rect 3593 -184 3613 -150
rect 3613 -184 3645 -150
rect 3657 -184 3685 -150
rect 3685 -184 3709 -150
rect 3721 -184 3757 -150
rect 3757 -184 3773 -150
rect 3785 -184 3791 -150
rect 3791 -184 3829 -150
rect 3829 -184 3837 -150
rect 3849 -184 3863 -150
rect 3863 -184 3901 -150
rect 3913 -184 3935 -150
rect 3935 -184 3965 -150
rect 3977 -184 4007 -150
rect 4007 -184 4029 -150
rect 3593 -194 3645 -184
rect 3657 -194 3709 -184
rect 3721 -194 3773 -184
rect 3785 -194 3837 -184
rect 3849 -194 3901 -184
rect 3913 -194 3965 -184
rect 3977 -194 4029 -184
rect 4041 -150 4093 -142
rect 4041 -184 4045 -150
rect 4045 -184 4079 -150
rect 4079 -184 4093 -150
rect 4041 -194 4093 -184
<< metal2 >>
rect 126 620 188 622
rect 318 620 380 622
rect 510 620 572 622
rect 702 620 764 622
rect 894 620 956 622
rect 1086 620 1148 622
rect 1278 620 1340 622
rect 1470 620 1532 622
rect 1662 620 1724 622
rect 1854 620 1916 622
rect 2046 620 2108 622
rect 2238 620 2300 622
rect 2430 620 2492 622
rect 2622 620 2684 622
rect 2814 620 2876 622
rect 3006 620 3068 622
rect 3198 620 3260 622
rect 3390 620 3452 622
rect 3582 620 3644 622
rect 3774 620 3836 622
rect 3966 620 4028 622
rect 126 611 190 620
rect 126 596 132 611
rect 184 596 190 611
rect 126 540 130 596
rect 186 540 190 596
rect 126 516 132 540
rect 184 516 190 540
rect 126 460 130 516
rect 186 460 190 516
rect 126 436 132 460
rect 184 436 190 460
rect 126 380 130 436
rect 186 380 190 436
rect 126 367 132 380
rect 184 367 190 380
rect 126 354 190 367
rect 318 611 382 620
rect 318 596 324 611
rect 376 596 382 611
rect 318 540 322 596
rect 378 540 382 596
rect 318 516 324 540
rect 376 516 382 540
rect 318 460 322 516
rect 378 460 382 516
rect 318 436 324 460
rect 376 436 382 460
rect 318 380 322 436
rect 378 380 382 436
rect 318 367 324 380
rect 376 367 382 380
rect 318 354 382 367
rect 510 611 574 620
rect 510 596 516 611
rect 568 596 574 611
rect 510 540 514 596
rect 570 540 574 596
rect 510 516 516 540
rect 568 516 574 540
rect 510 460 514 516
rect 570 460 574 516
rect 510 436 516 460
rect 568 436 574 460
rect 510 380 514 436
rect 570 380 574 436
rect 510 367 516 380
rect 568 367 574 380
rect 510 354 574 367
rect 702 611 766 620
rect 702 596 708 611
rect 760 596 766 611
rect 702 540 706 596
rect 762 540 766 596
rect 702 516 708 540
rect 760 516 766 540
rect 702 460 706 516
rect 762 460 766 516
rect 702 436 708 460
rect 760 436 766 460
rect 702 380 706 436
rect 762 380 766 436
rect 702 367 708 380
rect 760 367 766 380
rect 702 354 766 367
rect 894 611 958 620
rect 894 596 900 611
rect 952 596 958 611
rect 894 540 898 596
rect 954 540 958 596
rect 894 516 900 540
rect 952 516 958 540
rect 894 460 898 516
rect 954 460 958 516
rect 894 436 900 460
rect 952 436 958 460
rect 894 380 898 436
rect 954 380 958 436
rect 894 367 900 380
rect 952 367 958 380
rect 894 354 958 367
rect 1086 611 1150 620
rect 1086 596 1092 611
rect 1144 596 1150 611
rect 1086 540 1090 596
rect 1146 540 1150 596
rect 1086 516 1092 540
rect 1144 516 1150 540
rect 1086 460 1090 516
rect 1146 460 1150 516
rect 1086 436 1092 460
rect 1144 436 1150 460
rect 1086 380 1090 436
rect 1146 380 1150 436
rect 1086 367 1092 380
rect 1144 367 1150 380
rect 1086 354 1150 367
rect 1278 611 1342 620
rect 1278 596 1284 611
rect 1336 596 1342 611
rect 1278 540 1282 596
rect 1338 540 1342 596
rect 1278 516 1284 540
rect 1336 516 1342 540
rect 1278 460 1282 516
rect 1338 460 1342 516
rect 1278 436 1284 460
rect 1336 436 1342 460
rect 1278 380 1282 436
rect 1338 380 1342 436
rect 1278 367 1284 380
rect 1336 367 1342 380
rect 1278 354 1342 367
rect 1470 611 1534 620
rect 1470 596 1476 611
rect 1528 596 1534 611
rect 1470 540 1474 596
rect 1530 540 1534 596
rect 1470 516 1476 540
rect 1528 516 1534 540
rect 1470 460 1474 516
rect 1530 460 1534 516
rect 1470 436 1476 460
rect 1528 436 1534 460
rect 1470 380 1474 436
rect 1530 380 1534 436
rect 1470 367 1476 380
rect 1528 367 1534 380
rect 1470 354 1534 367
rect 1662 611 1726 620
rect 1662 596 1668 611
rect 1720 596 1726 611
rect 1662 540 1666 596
rect 1722 540 1726 596
rect 1662 516 1668 540
rect 1720 516 1726 540
rect 1662 460 1666 516
rect 1722 460 1726 516
rect 1662 436 1668 460
rect 1720 436 1726 460
rect 1662 380 1666 436
rect 1722 380 1726 436
rect 1662 367 1668 380
rect 1720 367 1726 380
rect 1662 354 1726 367
rect 1854 611 1918 620
rect 1854 596 1860 611
rect 1912 596 1918 611
rect 1854 540 1858 596
rect 1914 540 1918 596
rect 1854 516 1860 540
rect 1912 516 1918 540
rect 1854 460 1858 516
rect 1914 460 1918 516
rect 1854 436 1860 460
rect 1912 436 1918 460
rect 1854 380 1858 436
rect 1914 380 1918 436
rect 1854 367 1860 380
rect 1912 367 1918 380
rect 1854 354 1918 367
rect 2046 611 2110 620
rect 2046 596 2052 611
rect 2104 596 2110 611
rect 2046 540 2050 596
rect 2106 540 2110 596
rect 2046 516 2052 540
rect 2104 516 2110 540
rect 2046 460 2050 516
rect 2106 460 2110 516
rect 2046 436 2052 460
rect 2104 436 2110 460
rect 2046 380 2050 436
rect 2106 380 2110 436
rect 2046 367 2052 380
rect 2104 367 2110 380
rect 2046 354 2110 367
rect 2238 611 2302 620
rect 2238 596 2244 611
rect 2296 596 2302 611
rect 2238 540 2242 596
rect 2298 540 2302 596
rect 2238 516 2244 540
rect 2296 516 2302 540
rect 2238 460 2242 516
rect 2298 460 2302 516
rect 2238 436 2244 460
rect 2296 436 2302 460
rect 2238 380 2242 436
rect 2298 380 2302 436
rect 2238 367 2244 380
rect 2296 367 2302 380
rect 2238 354 2302 367
rect 2430 611 2494 620
rect 2430 596 2436 611
rect 2488 596 2494 611
rect 2430 540 2434 596
rect 2490 540 2494 596
rect 2430 516 2436 540
rect 2488 516 2494 540
rect 2430 460 2434 516
rect 2490 460 2494 516
rect 2430 436 2436 460
rect 2488 436 2494 460
rect 2430 380 2434 436
rect 2490 380 2494 436
rect 2430 367 2436 380
rect 2488 367 2494 380
rect 2430 354 2494 367
rect 2622 611 2686 620
rect 2622 596 2628 611
rect 2680 596 2686 611
rect 2622 540 2626 596
rect 2682 540 2686 596
rect 2622 516 2628 540
rect 2680 516 2686 540
rect 2622 460 2626 516
rect 2682 460 2686 516
rect 2622 436 2628 460
rect 2680 436 2686 460
rect 2622 380 2626 436
rect 2682 380 2686 436
rect 2622 367 2628 380
rect 2680 367 2686 380
rect 2622 354 2686 367
rect 2814 611 2878 620
rect 2814 596 2820 611
rect 2872 596 2878 611
rect 2814 540 2818 596
rect 2874 540 2878 596
rect 2814 516 2820 540
rect 2872 516 2878 540
rect 2814 460 2818 516
rect 2874 460 2878 516
rect 2814 436 2820 460
rect 2872 436 2878 460
rect 2814 380 2818 436
rect 2874 380 2878 436
rect 2814 367 2820 380
rect 2872 367 2878 380
rect 2814 354 2878 367
rect 3006 611 3070 620
rect 3006 596 3012 611
rect 3064 596 3070 611
rect 3006 540 3010 596
rect 3066 540 3070 596
rect 3006 516 3012 540
rect 3064 516 3070 540
rect 3006 460 3010 516
rect 3066 460 3070 516
rect 3006 436 3012 460
rect 3064 436 3070 460
rect 3006 380 3010 436
rect 3066 380 3070 436
rect 3006 367 3012 380
rect 3064 367 3070 380
rect 3006 354 3070 367
rect 3198 611 3262 620
rect 3198 596 3204 611
rect 3256 596 3262 611
rect 3198 540 3202 596
rect 3258 540 3262 596
rect 3198 516 3204 540
rect 3256 516 3262 540
rect 3198 460 3202 516
rect 3258 460 3262 516
rect 3198 436 3204 460
rect 3256 436 3262 460
rect 3198 380 3202 436
rect 3258 380 3262 436
rect 3198 367 3204 380
rect 3256 367 3262 380
rect 3198 354 3262 367
rect 3390 611 3454 620
rect 3390 596 3396 611
rect 3448 596 3454 611
rect 3390 540 3394 596
rect 3450 540 3454 596
rect 3390 516 3396 540
rect 3448 516 3454 540
rect 3390 460 3394 516
rect 3450 460 3454 516
rect 3390 436 3396 460
rect 3448 436 3454 460
rect 3390 380 3394 436
rect 3450 380 3454 436
rect 3390 367 3396 380
rect 3448 367 3454 380
rect 3390 354 3454 367
rect 3582 611 3646 620
rect 3582 596 3588 611
rect 3640 596 3646 611
rect 3582 540 3586 596
rect 3642 540 3646 596
rect 3582 516 3588 540
rect 3640 516 3646 540
rect 3582 460 3586 516
rect 3642 460 3646 516
rect 3582 436 3588 460
rect 3640 436 3646 460
rect 3582 380 3586 436
rect 3642 380 3646 436
rect 3582 367 3588 380
rect 3640 367 3646 380
rect 3582 354 3646 367
rect 3774 611 3838 620
rect 3774 596 3780 611
rect 3832 596 3838 611
rect 3774 540 3778 596
rect 3834 540 3838 596
rect 3774 516 3780 540
rect 3832 516 3838 540
rect 3774 460 3778 516
rect 3834 460 3838 516
rect 3774 436 3780 460
rect 3832 436 3838 460
rect 3774 380 3778 436
rect 3834 380 3838 436
rect 3774 367 3780 380
rect 3832 367 3838 380
rect 3774 354 3838 367
rect 3966 611 4030 620
rect 3966 596 3972 611
rect 4024 596 4030 611
rect 3966 540 3970 596
rect 4026 540 4030 596
rect 3966 516 3972 540
rect 4024 516 4030 540
rect 3966 460 3970 516
rect 4026 460 4030 516
rect 3966 436 3972 460
rect 4024 436 4030 460
rect 3966 380 3970 436
rect 4026 380 4030 436
rect 3966 367 3972 380
rect 4024 367 4030 380
rect 3966 354 4030 367
rect 30 279 94 284
rect 30 227 36 279
rect 88 227 94 279
rect 30 215 94 227
rect 30 163 36 215
rect 88 163 94 215
rect 30 151 94 163
rect 30 99 36 151
rect 88 99 94 151
rect 30 87 94 99
rect 30 35 36 87
rect 88 35 94 87
rect 30 -76 94 35
rect 222 279 286 284
rect 222 227 228 279
rect 280 227 286 279
rect 222 215 286 227
rect 222 163 228 215
rect 280 163 286 215
rect 222 151 286 163
rect 222 99 228 151
rect 280 99 286 151
rect 222 87 286 99
rect 222 35 228 87
rect 280 35 286 87
rect 222 -76 286 35
rect 414 279 478 284
rect 414 227 420 279
rect 472 227 478 279
rect 414 215 478 227
rect 414 163 420 215
rect 472 163 478 215
rect 414 151 478 163
rect 414 99 420 151
rect 472 99 478 151
rect 414 87 478 99
rect 414 35 420 87
rect 472 35 478 87
rect 414 -76 478 35
rect 606 279 670 284
rect 606 227 612 279
rect 664 227 670 279
rect 606 215 670 227
rect 606 163 612 215
rect 664 163 670 215
rect 606 151 670 163
rect 606 99 612 151
rect 664 99 670 151
rect 606 87 670 99
rect 606 35 612 87
rect 664 35 670 87
rect 606 -76 670 35
rect 798 279 862 284
rect 798 227 804 279
rect 856 227 862 279
rect 798 215 862 227
rect 798 163 804 215
rect 856 163 862 215
rect 798 151 862 163
rect 798 99 804 151
rect 856 99 862 151
rect 798 87 862 99
rect 798 35 804 87
rect 856 35 862 87
rect 798 -76 862 35
rect 990 279 1054 284
rect 990 227 996 279
rect 1048 227 1054 279
rect 990 215 1054 227
rect 990 163 996 215
rect 1048 163 1054 215
rect 990 151 1054 163
rect 990 99 996 151
rect 1048 99 1054 151
rect 990 87 1054 99
rect 990 35 996 87
rect 1048 35 1054 87
rect 990 -76 1054 35
rect 1182 279 1246 284
rect 1182 227 1188 279
rect 1240 227 1246 279
rect 1182 215 1246 227
rect 1182 163 1188 215
rect 1240 163 1246 215
rect 1182 151 1246 163
rect 1182 99 1188 151
rect 1240 99 1246 151
rect 1182 87 1246 99
rect 1182 35 1188 87
rect 1240 35 1246 87
rect 1182 -76 1246 35
rect 1374 279 1438 284
rect 1374 227 1380 279
rect 1432 227 1438 279
rect 1374 215 1438 227
rect 1374 163 1380 215
rect 1432 163 1438 215
rect 1374 151 1438 163
rect 1374 99 1380 151
rect 1432 99 1438 151
rect 1374 87 1438 99
rect 1374 35 1380 87
rect 1432 35 1438 87
rect 1374 -76 1438 35
rect 1566 279 1630 284
rect 1566 227 1572 279
rect 1624 227 1630 279
rect 1566 215 1630 227
rect 1566 163 1572 215
rect 1624 163 1630 215
rect 1566 151 1630 163
rect 1566 99 1572 151
rect 1624 99 1630 151
rect 1566 87 1630 99
rect 1566 35 1572 87
rect 1624 35 1630 87
rect 1566 -76 1630 35
rect 1758 279 1822 284
rect 1758 227 1764 279
rect 1816 227 1822 279
rect 1758 215 1822 227
rect 1758 163 1764 215
rect 1816 163 1822 215
rect 1758 151 1822 163
rect 1758 99 1764 151
rect 1816 99 1822 151
rect 1758 87 1822 99
rect 1758 35 1764 87
rect 1816 35 1822 87
rect 1758 -76 1822 35
rect 1950 279 2014 284
rect 1950 227 1956 279
rect 2008 227 2014 279
rect 1950 215 2014 227
rect 1950 163 1956 215
rect 2008 163 2014 215
rect 1950 151 2014 163
rect 1950 99 1956 151
rect 2008 99 2014 151
rect 1950 87 2014 99
rect 1950 35 1956 87
rect 2008 35 2014 87
rect 1950 -76 2014 35
rect 2142 279 2206 284
rect 2142 227 2148 279
rect 2200 227 2206 279
rect 2142 215 2206 227
rect 2142 163 2148 215
rect 2200 163 2206 215
rect 2142 151 2206 163
rect 2142 99 2148 151
rect 2200 99 2206 151
rect 2142 87 2206 99
rect 2142 35 2148 87
rect 2200 35 2206 87
rect 2142 -76 2206 35
rect 2334 279 2398 284
rect 2334 227 2340 279
rect 2392 227 2398 279
rect 2334 215 2398 227
rect 2334 163 2340 215
rect 2392 163 2398 215
rect 2334 151 2398 163
rect 2334 99 2340 151
rect 2392 99 2398 151
rect 2334 87 2398 99
rect 2334 35 2340 87
rect 2392 35 2398 87
rect 2334 -76 2398 35
rect 2526 279 2590 284
rect 2526 227 2532 279
rect 2584 227 2590 279
rect 2526 215 2590 227
rect 2526 163 2532 215
rect 2584 163 2590 215
rect 2526 151 2590 163
rect 2526 99 2532 151
rect 2584 99 2590 151
rect 2526 87 2590 99
rect 2526 35 2532 87
rect 2584 35 2590 87
rect 2526 -76 2590 35
rect 2718 279 2782 284
rect 2718 227 2724 279
rect 2776 227 2782 279
rect 2718 215 2782 227
rect 2718 163 2724 215
rect 2776 163 2782 215
rect 2718 151 2782 163
rect 2718 99 2724 151
rect 2776 99 2782 151
rect 2718 87 2782 99
rect 2718 35 2724 87
rect 2776 35 2782 87
rect 2718 -76 2782 35
rect 2910 279 2974 284
rect 2910 227 2916 279
rect 2968 227 2974 279
rect 2910 215 2974 227
rect 2910 163 2916 215
rect 2968 163 2974 215
rect 2910 151 2974 163
rect 2910 99 2916 151
rect 2968 99 2974 151
rect 2910 87 2974 99
rect 2910 35 2916 87
rect 2968 35 2974 87
rect 2910 -76 2974 35
rect 3102 279 3166 284
rect 3102 227 3108 279
rect 3160 227 3166 279
rect 3102 215 3166 227
rect 3102 163 3108 215
rect 3160 163 3166 215
rect 3102 151 3166 163
rect 3102 99 3108 151
rect 3160 99 3166 151
rect 3102 87 3166 99
rect 3102 35 3108 87
rect 3160 35 3166 87
rect 3102 -76 3166 35
rect 3294 279 3358 284
rect 3294 227 3300 279
rect 3352 227 3358 279
rect 3294 215 3358 227
rect 3294 163 3300 215
rect 3352 163 3358 215
rect 3294 151 3358 163
rect 3294 99 3300 151
rect 3352 99 3358 151
rect 3294 87 3358 99
rect 3294 35 3300 87
rect 3352 35 3358 87
rect 3294 -76 3358 35
rect 3486 279 3550 284
rect 3486 227 3492 279
rect 3544 227 3550 279
rect 3486 215 3550 227
rect 3486 163 3492 215
rect 3544 163 3550 215
rect 3486 151 3550 163
rect 3486 99 3492 151
rect 3544 99 3550 151
rect 3486 87 3550 99
rect 3486 35 3492 87
rect 3544 35 3550 87
rect 3486 -76 3550 35
rect 3678 279 3742 284
rect 3678 227 3684 279
rect 3736 227 3742 279
rect 3678 215 3742 227
rect 3678 163 3684 215
rect 3736 163 3742 215
rect 3678 151 3742 163
rect 3678 99 3684 151
rect 3736 99 3742 151
rect 3678 87 3742 99
rect 3678 35 3684 87
rect 3736 35 3742 87
rect 3678 -76 3742 35
rect 3870 279 3934 284
rect 3870 227 3876 279
rect 3928 227 3934 279
rect 3870 215 3934 227
rect 3870 163 3876 215
rect 3928 163 3934 215
rect 3870 151 3934 163
rect 3870 99 3876 151
rect 3928 99 3934 151
rect 3870 87 3934 99
rect 3870 35 3876 87
rect 3928 35 3934 87
rect 3870 -76 3934 35
rect 4062 279 4126 284
rect 4062 227 4068 279
rect 4120 227 4126 279
rect 4062 215 4126 227
rect 4062 163 4068 215
rect 4120 163 4126 215
rect 4062 151 4126 163
rect 4062 99 4068 151
rect 4120 99 4126 151
rect 4062 87 4126 99
rect 4062 35 4068 87
rect 4120 35 4126 87
rect 4062 -76 4126 35
rect 24 -142 4130 -76
rect 24 -194 73 -142
rect 125 -194 137 -142
rect 189 -194 201 -142
rect 253 -194 265 -142
rect 317 -194 329 -142
rect 381 -194 393 -142
rect 445 -194 457 -142
rect 509 -194 521 -142
rect 573 -194 585 -142
rect 637 -194 649 -142
rect 701 -194 713 -142
rect 765 -194 777 -142
rect 829 -194 841 -142
rect 893 -194 905 -142
rect 957 -194 969 -142
rect 1021 -194 1033 -142
rect 1085 -194 1097 -142
rect 1149 -194 1161 -142
rect 1213 -194 1225 -142
rect 1277 -194 1289 -142
rect 1341 -194 1353 -142
rect 1405 -194 1417 -142
rect 1469 -194 1481 -142
rect 1533 -194 1545 -142
rect 1597 -194 1609 -142
rect 1661 -194 1673 -142
rect 1725 -194 1737 -142
rect 1789 -194 1801 -142
rect 1853 -194 1865 -142
rect 1917 -194 1929 -142
rect 1981 -194 1993 -142
rect 2045 -194 2057 -142
rect 2109 -194 2121 -142
rect 2173 -194 2185 -142
rect 2237 -194 2249 -142
rect 2301 -194 2313 -142
rect 2365 -194 2377 -142
rect 2429 -194 2441 -142
rect 2493 -194 2505 -142
rect 2557 -194 2569 -142
rect 2621 -194 2633 -142
rect 2685 -194 2697 -142
rect 2749 -194 2761 -142
rect 2813 -194 2825 -142
rect 2877 -194 2889 -142
rect 2941 -194 2953 -142
rect 3005 -194 3017 -142
rect 3069 -194 3081 -142
rect 3133 -194 3145 -142
rect 3197 -194 3209 -142
rect 3261 -194 3273 -142
rect 3325 -194 3337 -142
rect 3389 -194 3401 -142
rect 3453 -194 3465 -142
rect 3517 -194 3529 -142
rect 3581 -194 3593 -142
rect 3645 -194 3657 -142
rect 3709 -194 3721 -142
rect 3773 -194 3785 -142
rect 3837 -194 3849 -142
rect 3901 -194 3913 -142
rect 3965 -194 3977 -142
rect 4029 -194 4041 -142
rect 4093 -194 4130 -142
rect 24 -284 4130 -194
rect 24 -320 4128 -284
<< via2 >>
rect 130 559 132 596
rect 132 559 184 596
rect 184 559 186 596
rect 130 547 186 559
rect 130 540 132 547
rect 132 540 184 547
rect 184 540 186 547
rect 130 495 132 516
rect 132 495 184 516
rect 184 495 186 516
rect 130 483 186 495
rect 130 460 132 483
rect 132 460 184 483
rect 184 460 186 483
rect 130 431 132 436
rect 132 431 184 436
rect 184 431 186 436
rect 130 419 186 431
rect 130 380 132 419
rect 132 380 184 419
rect 184 380 186 419
rect 322 559 324 596
rect 324 559 376 596
rect 376 559 378 596
rect 322 547 378 559
rect 322 540 324 547
rect 324 540 376 547
rect 376 540 378 547
rect 322 495 324 516
rect 324 495 376 516
rect 376 495 378 516
rect 322 483 378 495
rect 322 460 324 483
rect 324 460 376 483
rect 376 460 378 483
rect 322 431 324 436
rect 324 431 376 436
rect 376 431 378 436
rect 322 419 378 431
rect 322 380 324 419
rect 324 380 376 419
rect 376 380 378 419
rect 514 559 516 596
rect 516 559 568 596
rect 568 559 570 596
rect 514 547 570 559
rect 514 540 516 547
rect 516 540 568 547
rect 568 540 570 547
rect 514 495 516 516
rect 516 495 568 516
rect 568 495 570 516
rect 514 483 570 495
rect 514 460 516 483
rect 516 460 568 483
rect 568 460 570 483
rect 514 431 516 436
rect 516 431 568 436
rect 568 431 570 436
rect 514 419 570 431
rect 514 380 516 419
rect 516 380 568 419
rect 568 380 570 419
rect 706 559 708 596
rect 708 559 760 596
rect 760 559 762 596
rect 706 547 762 559
rect 706 540 708 547
rect 708 540 760 547
rect 760 540 762 547
rect 706 495 708 516
rect 708 495 760 516
rect 760 495 762 516
rect 706 483 762 495
rect 706 460 708 483
rect 708 460 760 483
rect 760 460 762 483
rect 706 431 708 436
rect 708 431 760 436
rect 760 431 762 436
rect 706 419 762 431
rect 706 380 708 419
rect 708 380 760 419
rect 760 380 762 419
rect 898 559 900 596
rect 900 559 952 596
rect 952 559 954 596
rect 898 547 954 559
rect 898 540 900 547
rect 900 540 952 547
rect 952 540 954 547
rect 898 495 900 516
rect 900 495 952 516
rect 952 495 954 516
rect 898 483 954 495
rect 898 460 900 483
rect 900 460 952 483
rect 952 460 954 483
rect 898 431 900 436
rect 900 431 952 436
rect 952 431 954 436
rect 898 419 954 431
rect 898 380 900 419
rect 900 380 952 419
rect 952 380 954 419
rect 1090 559 1092 596
rect 1092 559 1144 596
rect 1144 559 1146 596
rect 1090 547 1146 559
rect 1090 540 1092 547
rect 1092 540 1144 547
rect 1144 540 1146 547
rect 1090 495 1092 516
rect 1092 495 1144 516
rect 1144 495 1146 516
rect 1090 483 1146 495
rect 1090 460 1092 483
rect 1092 460 1144 483
rect 1144 460 1146 483
rect 1090 431 1092 436
rect 1092 431 1144 436
rect 1144 431 1146 436
rect 1090 419 1146 431
rect 1090 380 1092 419
rect 1092 380 1144 419
rect 1144 380 1146 419
rect 1282 559 1284 596
rect 1284 559 1336 596
rect 1336 559 1338 596
rect 1282 547 1338 559
rect 1282 540 1284 547
rect 1284 540 1336 547
rect 1336 540 1338 547
rect 1282 495 1284 516
rect 1284 495 1336 516
rect 1336 495 1338 516
rect 1282 483 1338 495
rect 1282 460 1284 483
rect 1284 460 1336 483
rect 1336 460 1338 483
rect 1282 431 1284 436
rect 1284 431 1336 436
rect 1336 431 1338 436
rect 1282 419 1338 431
rect 1282 380 1284 419
rect 1284 380 1336 419
rect 1336 380 1338 419
rect 1474 559 1476 596
rect 1476 559 1528 596
rect 1528 559 1530 596
rect 1474 547 1530 559
rect 1474 540 1476 547
rect 1476 540 1528 547
rect 1528 540 1530 547
rect 1474 495 1476 516
rect 1476 495 1528 516
rect 1528 495 1530 516
rect 1474 483 1530 495
rect 1474 460 1476 483
rect 1476 460 1528 483
rect 1528 460 1530 483
rect 1474 431 1476 436
rect 1476 431 1528 436
rect 1528 431 1530 436
rect 1474 419 1530 431
rect 1474 380 1476 419
rect 1476 380 1528 419
rect 1528 380 1530 419
rect 1666 559 1668 596
rect 1668 559 1720 596
rect 1720 559 1722 596
rect 1666 547 1722 559
rect 1666 540 1668 547
rect 1668 540 1720 547
rect 1720 540 1722 547
rect 1666 495 1668 516
rect 1668 495 1720 516
rect 1720 495 1722 516
rect 1666 483 1722 495
rect 1666 460 1668 483
rect 1668 460 1720 483
rect 1720 460 1722 483
rect 1666 431 1668 436
rect 1668 431 1720 436
rect 1720 431 1722 436
rect 1666 419 1722 431
rect 1666 380 1668 419
rect 1668 380 1720 419
rect 1720 380 1722 419
rect 1858 559 1860 596
rect 1860 559 1912 596
rect 1912 559 1914 596
rect 1858 547 1914 559
rect 1858 540 1860 547
rect 1860 540 1912 547
rect 1912 540 1914 547
rect 1858 495 1860 516
rect 1860 495 1912 516
rect 1912 495 1914 516
rect 1858 483 1914 495
rect 1858 460 1860 483
rect 1860 460 1912 483
rect 1912 460 1914 483
rect 1858 431 1860 436
rect 1860 431 1912 436
rect 1912 431 1914 436
rect 1858 419 1914 431
rect 1858 380 1860 419
rect 1860 380 1912 419
rect 1912 380 1914 419
rect 2050 559 2052 596
rect 2052 559 2104 596
rect 2104 559 2106 596
rect 2050 547 2106 559
rect 2050 540 2052 547
rect 2052 540 2104 547
rect 2104 540 2106 547
rect 2050 495 2052 516
rect 2052 495 2104 516
rect 2104 495 2106 516
rect 2050 483 2106 495
rect 2050 460 2052 483
rect 2052 460 2104 483
rect 2104 460 2106 483
rect 2050 431 2052 436
rect 2052 431 2104 436
rect 2104 431 2106 436
rect 2050 419 2106 431
rect 2050 380 2052 419
rect 2052 380 2104 419
rect 2104 380 2106 419
rect 2242 559 2244 596
rect 2244 559 2296 596
rect 2296 559 2298 596
rect 2242 547 2298 559
rect 2242 540 2244 547
rect 2244 540 2296 547
rect 2296 540 2298 547
rect 2242 495 2244 516
rect 2244 495 2296 516
rect 2296 495 2298 516
rect 2242 483 2298 495
rect 2242 460 2244 483
rect 2244 460 2296 483
rect 2296 460 2298 483
rect 2242 431 2244 436
rect 2244 431 2296 436
rect 2296 431 2298 436
rect 2242 419 2298 431
rect 2242 380 2244 419
rect 2244 380 2296 419
rect 2296 380 2298 419
rect 2434 559 2436 596
rect 2436 559 2488 596
rect 2488 559 2490 596
rect 2434 547 2490 559
rect 2434 540 2436 547
rect 2436 540 2488 547
rect 2488 540 2490 547
rect 2434 495 2436 516
rect 2436 495 2488 516
rect 2488 495 2490 516
rect 2434 483 2490 495
rect 2434 460 2436 483
rect 2436 460 2488 483
rect 2488 460 2490 483
rect 2434 431 2436 436
rect 2436 431 2488 436
rect 2488 431 2490 436
rect 2434 419 2490 431
rect 2434 380 2436 419
rect 2436 380 2488 419
rect 2488 380 2490 419
rect 2626 559 2628 596
rect 2628 559 2680 596
rect 2680 559 2682 596
rect 2626 547 2682 559
rect 2626 540 2628 547
rect 2628 540 2680 547
rect 2680 540 2682 547
rect 2626 495 2628 516
rect 2628 495 2680 516
rect 2680 495 2682 516
rect 2626 483 2682 495
rect 2626 460 2628 483
rect 2628 460 2680 483
rect 2680 460 2682 483
rect 2626 431 2628 436
rect 2628 431 2680 436
rect 2680 431 2682 436
rect 2626 419 2682 431
rect 2626 380 2628 419
rect 2628 380 2680 419
rect 2680 380 2682 419
rect 2818 559 2820 596
rect 2820 559 2872 596
rect 2872 559 2874 596
rect 2818 547 2874 559
rect 2818 540 2820 547
rect 2820 540 2872 547
rect 2872 540 2874 547
rect 2818 495 2820 516
rect 2820 495 2872 516
rect 2872 495 2874 516
rect 2818 483 2874 495
rect 2818 460 2820 483
rect 2820 460 2872 483
rect 2872 460 2874 483
rect 2818 431 2820 436
rect 2820 431 2872 436
rect 2872 431 2874 436
rect 2818 419 2874 431
rect 2818 380 2820 419
rect 2820 380 2872 419
rect 2872 380 2874 419
rect 3010 559 3012 596
rect 3012 559 3064 596
rect 3064 559 3066 596
rect 3010 547 3066 559
rect 3010 540 3012 547
rect 3012 540 3064 547
rect 3064 540 3066 547
rect 3010 495 3012 516
rect 3012 495 3064 516
rect 3064 495 3066 516
rect 3010 483 3066 495
rect 3010 460 3012 483
rect 3012 460 3064 483
rect 3064 460 3066 483
rect 3010 431 3012 436
rect 3012 431 3064 436
rect 3064 431 3066 436
rect 3010 419 3066 431
rect 3010 380 3012 419
rect 3012 380 3064 419
rect 3064 380 3066 419
rect 3202 559 3204 596
rect 3204 559 3256 596
rect 3256 559 3258 596
rect 3202 547 3258 559
rect 3202 540 3204 547
rect 3204 540 3256 547
rect 3256 540 3258 547
rect 3202 495 3204 516
rect 3204 495 3256 516
rect 3256 495 3258 516
rect 3202 483 3258 495
rect 3202 460 3204 483
rect 3204 460 3256 483
rect 3256 460 3258 483
rect 3202 431 3204 436
rect 3204 431 3256 436
rect 3256 431 3258 436
rect 3202 419 3258 431
rect 3202 380 3204 419
rect 3204 380 3256 419
rect 3256 380 3258 419
rect 3394 559 3396 596
rect 3396 559 3448 596
rect 3448 559 3450 596
rect 3394 547 3450 559
rect 3394 540 3396 547
rect 3396 540 3448 547
rect 3448 540 3450 547
rect 3394 495 3396 516
rect 3396 495 3448 516
rect 3448 495 3450 516
rect 3394 483 3450 495
rect 3394 460 3396 483
rect 3396 460 3448 483
rect 3448 460 3450 483
rect 3394 431 3396 436
rect 3396 431 3448 436
rect 3448 431 3450 436
rect 3394 419 3450 431
rect 3394 380 3396 419
rect 3396 380 3448 419
rect 3448 380 3450 419
rect 3586 559 3588 596
rect 3588 559 3640 596
rect 3640 559 3642 596
rect 3586 547 3642 559
rect 3586 540 3588 547
rect 3588 540 3640 547
rect 3640 540 3642 547
rect 3586 495 3588 516
rect 3588 495 3640 516
rect 3640 495 3642 516
rect 3586 483 3642 495
rect 3586 460 3588 483
rect 3588 460 3640 483
rect 3640 460 3642 483
rect 3586 431 3588 436
rect 3588 431 3640 436
rect 3640 431 3642 436
rect 3586 419 3642 431
rect 3586 380 3588 419
rect 3588 380 3640 419
rect 3640 380 3642 419
rect 3778 559 3780 596
rect 3780 559 3832 596
rect 3832 559 3834 596
rect 3778 547 3834 559
rect 3778 540 3780 547
rect 3780 540 3832 547
rect 3832 540 3834 547
rect 3778 495 3780 516
rect 3780 495 3832 516
rect 3832 495 3834 516
rect 3778 483 3834 495
rect 3778 460 3780 483
rect 3780 460 3832 483
rect 3832 460 3834 483
rect 3778 431 3780 436
rect 3780 431 3832 436
rect 3832 431 3834 436
rect 3778 419 3834 431
rect 3778 380 3780 419
rect 3780 380 3832 419
rect 3832 380 3834 419
rect 3970 559 3972 596
rect 3972 559 4024 596
rect 4024 559 4026 596
rect 3970 547 4026 559
rect 3970 540 3972 547
rect 3972 540 4024 547
rect 4024 540 4026 547
rect 3970 495 3972 516
rect 3972 495 4024 516
rect 4024 495 4026 516
rect 3970 483 4026 495
rect 3970 460 3972 483
rect 3972 460 4024 483
rect 4024 460 4026 483
rect 3970 431 3972 436
rect 3972 431 4024 436
rect 4024 431 4026 436
rect 3970 419 4026 431
rect 3970 380 3972 419
rect 3972 380 4024 419
rect 4024 380 4026 419
<< metal3 >>
rect 124 728 4032 814
rect 124 596 192 728
rect 124 540 130 596
rect 186 540 192 596
rect 124 516 192 540
rect 124 460 130 516
rect 186 460 192 516
rect 124 436 192 460
rect 124 380 130 436
rect 186 380 192 436
rect 124 354 192 380
rect 316 596 384 728
rect 316 540 322 596
rect 378 540 384 596
rect 316 516 384 540
rect 316 460 322 516
rect 378 460 384 516
rect 316 436 384 460
rect 316 380 322 436
rect 378 380 384 436
rect 316 354 384 380
rect 508 596 576 728
rect 508 540 514 596
rect 570 540 576 596
rect 508 516 576 540
rect 508 460 514 516
rect 570 460 576 516
rect 508 436 576 460
rect 508 380 514 436
rect 570 380 576 436
rect 508 354 576 380
rect 700 596 768 728
rect 700 540 706 596
rect 762 540 768 596
rect 700 516 768 540
rect 700 460 706 516
rect 762 460 768 516
rect 700 436 768 460
rect 700 380 706 436
rect 762 380 768 436
rect 700 354 768 380
rect 892 596 960 728
rect 892 540 898 596
rect 954 540 960 596
rect 892 516 960 540
rect 892 460 898 516
rect 954 460 960 516
rect 892 436 960 460
rect 892 380 898 436
rect 954 380 960 436
rect 892 354 960 380
rect 1084 596 1152 728
rect 1084 540 1090 596
rect 1146 540 1152 596
rect 1084 516 1152 540
rect 1084 460 1090 516
rect 1146 460 1152 516
rect 1084 436 1152 460
rect 1084 380 1090 436
rect 1146 380 1152 436
rect 1084 354 1152 380
rect 1276 596 1344 728
rect 1276 540 1282 596
rect 1338 540 1344 596
rect 1276 516 1344 540
rect 1276 460 1282 516
rect 1338 460 1344 516
rect 1276 436 1344 460
rect 1276 380 1282 436
rect 1338 380 1344 436
rect 1276 354 1344 380
rect 1468 596 1536 728
rect 1468 540 1474 596
rect 1530 540 1536 596
rect 1468 516 1536 540
rect 1468 460 1474 516
rect 1530 460 1536 516
rect 1468 436 1536 460
rect 1468 380 1474 436
rect 1530 380 1536 436
rect 1468 354 1536 380
rect 1660 596 1728 728
rect 1660 540 1666 596
rect 1722 540 1728 596
rect 1660 516 1728 540
rect 1660 460 1666 516
rect 1722 460 1728 516
rect 1660 436 1728 460
rect 1660 380 1666 436
rect 1722 380 1728 436
rect 1660 354 1728 380
rect 1852 596 1920 728
rect 1852 540 1858 596
rect 1914 540 1920 596
rect 1852 516 1920 540
rect 1852 460 1858 516
rect 1914 460 1920 516
rect 1852 436 1920 460
rect 1852 380 1858 436
rect 1914 380 1920 436
rect 1852 354 1920 380
rect 2044 596 2112 728
rect 2044 540 2050 596
rect 2106 540 2112 596
rect 2044 516 2112 540
rect 2044 460 2050 516
rect 2106 460 2112 516
rect 2044 436 2112 460
rect 2044 380 2050 436
rect 2106 380 2112 436
rect 2044 354 2112 380
rect 2236 596 2304 728
rect 2236 540 2242 596
rect 2298 540 2304 596
rect 2236 516 2304 540
rect 2236 460 2242 516
rect 2298 460 2304 516
rect 2236 436 2304 460
rect 2236 380 2242 436
rect 2298 380 2304 436
rect 2236 354 2304 380
rect 2428 596 2496 728
rect 2428 540 2434 596
rect 2490 540 2496 596
rect 2428 516 2496 540
rect 2428 460 2434 516
rect 2490 460 2496 516
rect 2428 436 2496 460
rect 2428 380 2434 436
rect 2490 380 2496 436
rect 2428 354 2496 380
rect 2620 596 2688 728
rect 2620 540 2626 596
rect 2682 540 2688 596
rect 2620 516 2688 540
rect 2620 460 2626 516
rect 2682 460 2688 516
rect 2620 436 2688 460
rect 2620 380 2626 436
rect 2682 380 2688 436
rect 2620 354 2688 380
rect 2812 596 2880 728
rect 2812 540 2818 596
rect 2874 540 2880 596
rect 2812 516 2880 540
rect 2812 460 2818 516
rect 2874 460 2880 516
rect 2812 436 2880 460
rect 2812 380 2818 436
rect 2874 380 2880 436
rect 2812 354 2880 380
rect 3004 596 3072 728
rect 3004 540 3010 596
rect 3066 540 3072 596
rect 3004 516 3072 540
rect 3004 460 3010 516
rect 3066 460 3072 516
rect 3004 436 3072 460
rect 3004 380 3010 436
rect 3066 380 3072 436
rect 3004 354 3072 380
rect 3196 596 3264 728
rect 3196 540 3202 596
rect 3258 540 3264 596
rect 3196 516 3264 540
rect 3196 460 3202 516
rect 3258 460 3264 516
rect 3196 436 3264 460
rect 3196 380 3202 436
rect 3258 380 3264 436
rect 3196 354 3264 380
rect 3388 596 3456 728
rect 3388 540 3394 596
rect 3450 540 3456 596
rect 3388 516 3456 540
rect 3388 460 3394 516
rect 3450 460 3456 516
rect 3388 436 3456 460
rect 3388 380 3394 436
rect 3450 380 3456 436
rect 3388 354 3456 380
rect 3580 596 3648 728
rect 3580 540 3586 596
rect 3642 540 3648 596
rect 3580 516 3648 540
rect 3580 460 3586 516
rect 3642 460 3648 516
rect 3580 436 3648 460
rect 3580 380 3586 436
rect 3642 380 3648 436
rect 3580 354 3648 380
rect 3772 596 3840 728
rect 3772 540 3778 596
rect 3834 540 3840 596
rect 3772 516 3840 540
rect 3772 460 3778 516
rect 3834 460 3840 516
rect 3772 436 3840 460
rect 3772 380 3778 436
rect 3834 380 3840 436
rect 3772 354 3840 380
rect 3964 596 4032 728
rect 3964 540 3970 596
rect 4026 540 4032 596
rect 3964 516 4032 540
rect 3964 460 3970 516
rect 4026 460 4032 516
rect 3964 436 4032 460
rect 3964 380 3970 436
rect 4026 380 4032 436
rect 3964 354 4032 380
use sky130_fd_pr__nfet_01v8_4PXCG5  sky130_fd_pr__nfet_01v8_4PXCG5_0
timestamp 1627926120
transform 1 0 2077 0 -1 323
box -2147 -474 2147 474
<< labels >>
rlabel metal2 s 28 -318 4124 -206 4 GND
port 1 nsew
rlabel metal1 s 80 656 3976 704 4 gate
port 2 nsew
rlabel metal3 s 124 748 4024 810 4 vl
port 3 nsew
<< end >>
