magic
tech sky130A
magscale 1 2
timestamp 1627036492
<< pwell >>
rect -3222 -1286 3222 1286
<< psubdiff >>
rect -3186 1216 3186 1250
rect -3186 -1216 -3152 1216
rect 3152 -1216 3186 1216
rect -3186 -1250 -3090 -1216
rect 3090 -1250 3186 -1216
<< psubdiffcont >>
rect -3090 -1250 3090 -1216
<< xpolycontact >>
rect -3056 688 -2986 1120
rect -3056 -1120 -2986 -688
rect -2738 688 -2668 1120
rect -2738 -1120 -2668 -688
rect -2420 688 -2350 1120
rect -2420 -1120 -2350 -688
rect -2102 688 -2032 1120
rect -2102 -1120 -2032 -688
rect -1784 688 -1714 1120
rect -1784 -1120 -1714 -688
rect -1466 688 -1396 1120
rect -1466 -1120 -1396 -688
rect -1148 688 -1078 1120
rect -1148 -1120 -1078 -688
rect -830 688 -760 1120
rect -830 -1120 -760 -688
rect -512 688 -442 1120
rect -512 -1120 -442 -688
rect -194 688 -124 1120
rect -194 -1120 -124 -688
rect 124 688 194 1120
rect 124 -1120 194 -688
rect 442 688 512 1120
rect 442 -1120 512 -688
rect 760 688 830 1120
rect 760 -1120 830 -688
rect 1078 688 1148 1120
rect 1078 -1120 1148 -688
rect 1396 688 1466 1120
rect 1396 -1120 1466 -688
rect 1714 688 1784 1120
rect 1714 -1120 1784 -688
rect 2032 688 2102 1120
rect 2032 -1120 2102 -688
rect 2350 688 2420 1120
rect 2350 -1120 2420 -688
rect 2668 688 2738 1120
rect 2668 -1120 2738 -688
rect 2986 688 3056 1120
rect 2986 -1120 3056 -688
<< xpolyres >>
rect -3056 -688 -2986 688
rect -2738 -688 -2668 688
rect -2420 -688 -2350 688
rect -2102 -688 -2032 688
rect -1784 -688 -1714 688
rect -1466 -688 -1396 688
rect -1148 -688 -1078 688
rect -830 -688 -760 688
rect -512 -688 -442 688
rect -194 -688 -124 688
rect 124 -688 194 688
rect 442 -688 512 688
rect 760 -688 830 688
rect 1078 -688 1148 688
rect 1396 -688 1466 688
rect 1714 -688 1784 688
rect 2032 -688 2102 688
rect 2350 -688 2420 688
rect 2668 -688 2738 688
rect 2986 -688 3056 688
<< locali >>
rect -3186 1216 3186 1250
rect -3186 -1216 -3152 1216
rect 3152 -1216 3186 1216
rect -3186 -1250 -3090 -1216
rect 3090 -1250 3186 -1216
<< viali >>
rect -3040 705 -3002 1102
rect -2722 705 -2684 1102
rect -2404 705 -2366 1102
rect -2086 705 -2048 1102
rect -1768 705 -1730 1102
rect -1450 705 -1412 1102
rect -1132 705 -1094 1102
rect -814 705 -776 1102
rect -496 705 -458 1102
rect -178 705 -140 1102
rect 140 705 178 1102
rect 458 705 496 1102
rect 776 705 814 1102
rect 1094 705 1132 1102
rect 1412 705 1450 1102
rect 1730 705 1768 1102
rect 2048 705 2086 1102
rect 2366 705 2404 1102
rect 2684 705 2722 1102
rect 3002 705 3040 1102
rect -3040 -1102 -3002 -705
rect -2722 -1102 -2684 -705
rect -2404 -1102 -2366 -705
rect -2086 -1102 -2048 -705
rect -1768 -1102 -1730 -705
rect -1450 -1102 -1412 -705
rect -1132 -1102 -1094 -705
rect -814 -1102 -776 -705
rect -496 -1102 -458 -705
rect -178 -1102 -140 -705
rect 140 -1102 178 -705
rect 458 -1102 496 -705
rect 776 -1102 814 -705
rect 1094 -1102 1132 -705
rect 1412 -1102 1450 -705
rect 1730 -1102 1768 -705
rect 2048 -1102 2086 -705
rect 2366 -1102 2404 -705
rect 2684 -1102 2722 -705
rect 3002 -1102 3040 -705
<< metal1 >>
rect -3046 1102 -2996 1114
rect -3046 705 -3040 1102
rect -3002 705 -2996 1102
rect -3046 693 -2996 705
rect -2728 1102 -2678 1114
rect -2728 705 -2722 1102
rect -2684 705 -2678 1102
rect -2728 693 -2678 705
rect -2410 1102 -2360 1114
rect -2410 705 -2404 1102
rect -2366 705 -2360 1102
rect -2410 693 -2360 705
rect -2092 1102 -2042 1114
rect -2092 705 -2086 1102
rect -2048 705 -2042 1102
rect -2092 693 -2042 705
rect -1774 1102 -1724 1114
rect -1774 705 -1768 1102
rect -1730 705 -1724 1102
rect -1774 693 -1724 705
rect -1456 1102 -1406 1114
rect -1456 705 -1450 1102
rect -1412 705 -1406 1102
rect -1456 693 -1406 705
rect -1138 1102 -1088 1114
rect -1138 705 -1132 1102
rect -1094 705 -1088 1102
rect -1138 693 -1088 705
rect -820 1102 -770 1114
rect -820 705 -814 1102
rect -776 705 -770 1102
rect -820 693 -770 705
rect -502 1102 -452 1114
rect -502 705 -496 1102
rect -458 705 -452 1102
rect -502 693 -452 705
rect -184 1102 -134 1114
rect -184 705 -178 1102
rect -140 705 -134 1102
rect -184 693 -134 705
rect 134 1102 184 1114
rect 134 705 140 1102
rect 178 705 184 1102
rect 134 693 184 705
rect 452 1102 502 1114
rect 452 705 458 1102
rect 496 705 502 1102
rect 452 693 502 705
rect 770 1102 820 1114
rect 770 705 776 1102
rect 814 705 820 1102
rect 770 693 820 705
rect 1088 1102 1138 1114
rect 1088 705 1094 1102
rect 1132 705 1138 1102
rect 1088 693 1138 705
rect 1406 1102 1456 1114
rect 1406 705 1412 1102
rect 1450 705 1456 1102
rect 1406 693 1456 705
rect 1724 1102 1774 1114
rect 1724 705 1730 1102
rect 1768 705 1774 1102
rect 1724 693 1774 705
rect 2042 1102 2092 1114
rect 2042 705 2048 1102
rect 2086 705 2092 1102
rect 2042 693 2092 705
rect 2360 1102 2410 1114
rect 2360 705 2366 1102
rect 2404 705 2410 1102
rect 2360 693 2410 705
rect 2678 1102 2728 1114
rect 2678 705 2684 1102
rect 2722 705 2728 1102
rect 2678 693 2728 705
rect 2996 1102 3046 1114
rect 2996 705 3002 1102
rect 3040 705 3046 1102
rect 2996 693 3046 705
rect -3046 -705 -2996 -693
rect -3046 -1102 -3040 -705
rect -3002 -1102 -2996 -705
rect -3046 -1114 -2996 -1102
rect -2728 -705 -2678 -693
rect -2728 -1102 -2722 -705
rect -2684 -1102 -2678 -705
rect -2728 -1114 -2678 -1102
rect -2410 -705 -2360 -693
rect -2410 -1102 -2404 -705
rect -2366 -1102 -2360 -705
rect -2410 -1114 -2360 -1102
rect -2092 -705 -2042 -693
rect -2092 -1102 -2086 -705
rect -2048 -1102 -2042 -705
rect -2092 -1114 -2042 -1102
rect -1774 -705 -1724 -693
rect -1774 -1102 -1768 -705
rect -1730 -1102 -1724 -705
rect -1774 -1114 -1724 -1102
rect -1456 -705 -1406 -693
rect -1456 -1102 -1450 -705
rect -1412 -1102 -1406 -705
rect -1456 -1114 -1406 -1102
rect -1138 -705 -1088 -693
rect -1138 -1102 -1132 -705
rect -1094 -1102 -1088 -705
rect -1138 -1114 -1088 -1102
rect -820 -705 -770 -693
rect -820 -1102 -814 -705
rect -776 -1102 -770 -705
rect -820 -1114 -770 -1102
rect -502 -705 -452 -693
rect -502 -1102 -496 -705
rect -458 -1102 -452 -705
rect -502 -1114 -452 -1102
rect -184 -705 -134 -693
rect -184 -1102 -178 -705
rect -140 -1102 -134 -705
rect -184 -1114 -134 -1102
rect 134 -705 184 -693
rect 134 -1102 140 -705
rect 178 -1102 184 -705
rect 134 -1114 184 -1102
rect 452 -705 502 -693
rect 452 -1102 458 -705
rect 496 -1102 502 -705
rect 452 -1114 502 -1102
rect 770 -705 820 -693
rect 770 -1102 776 -705
rect 814 -1102 820 -705
rect 770 -1114 820 -1102
rect 1088 -705 1138 -693
rect 1088 -1102 1094 -705
rect 1132 -1102 1138 -705
rect 1088 -1114 1138 -1102
rect 1406 -705 1456 -693
rect 1406 -1102 1412 -705
rect 1450 -1102 1456 -705
rect 1406 -1114 1456 -1102
rect 1724 -705 1774 -693
rect 1724 -1102 1730 -705
rect 1768 -1102 1774 -705
rect 1724 -1114 1774 -1102
rect 2042 -705 2092 -693
rect 2042 -1102 2048 -705
rect 2086 -1102 2092 -705
rect 2042 -1114 2092 -1102
rect 2360 -705 2410 -693
rect 2360 -1102 2366 -705
rect 2404 -1102 2410 -705
rect 2360 -1114 2410 -1102
rect 2678 -705 2728 -693
rect 2678 -1102 2684 -705
rect 2722 -1102 2728 -705
rect 2678 -1114 2728 -1102
rect 2996 -705 3046 -693
rect 2996 -1102 3002 -705
rect 3040 -1102 3046 -705
rect 2996 -1114 3046 -1102
<< res0p35 >>
rect -3058 -690 -2984 690
rect -2740 -690 -2666 690
rect -2422 -690 -2348 690
rect -2104 -690 -2030 690
rect -1786 -690 -1712 690
rect -1468 -690 -1394 690
rect -1150 -690 -1076 690
rect -832 -690 -758 690
rect -514 -690 -440 690
rect -196 -690 -122 690
rect 122 -690 196 690
rect 440 -690 514 690
rect 758 -690 832 690
rect 1076 -690 1150 690
rect 1394 -690 1468 690
rect 1712 -690 1786 690
rect 2030 -690 2104 690
rect 2348 -690 2422 690
rect 2666 -690 2740 690
rect 2984 -690 3058 690
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string FIXED_BBOX -3169 -1233 3169 1233
string parameters w 0.350 l 6.88 m 1 nx 20 wmin 0.350 lmin 0.50 rho 2000 val 40.0k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 0 grc 0 gtc 0 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
