magic
tech sky130A
magscale 1 2
timestamp 1627922418
<< xpolycontact >>
rect -35 343 35 775
rect -35 -775 35 -343
<< xpolyres >>
rect -35 -343 35 343
<< viali >>
rect -19 360 19 757
rect -19 -757 19 -360
<< metal1 >>
rect -25 757 25 769
rect -25 360 -19 757
rect 19 360 25 757
rect -25 348 25 360
rect -25 -360 25 -348
rect -25 -757 -19 -360
rect 19 -757 25 -360
rect -25 -769 25 -757
<< res0p35 >>
rect -37 -345 37 345
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 3.43 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 20.285k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
