magic
tech sky130A
magscale 1 2
timestamp 1626782926
<< error_p >>
rect -29 3671 29 3677
rect -29 3637 -17 3671
rect -29 3631 29 3637
rect -29 2543 29 2549
rect -29 2509 -17 2543
rect -29 2503 29 2509
rect -29 2435 29 2441
rect -29 2401 -17 2435
rect -29 2395 29 2401
rect -29 1307 29 1313
rect -29 1273 -17 1307
rect -29 1267 29 1273
rect -29 1199 29 1205
rect -29 1165 -17 1199
rect -29 1159 29 1165
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -1165 29 -1159
rect -29 -1199 -17 -1165
rect -29 -1205 29 -1199
rect -29 -1273 29 -1267
rect -29 -1307 -17 -1273
rect -29 -1313 29 -1307
rect -29 -2401 29 -2395
rect -29 -2435 -17 -2401
rect -29 -2441 29 -2435
rect -29 -2509 29 -2503
rect -29 -2543 -17 -2509
rect -29 -2549 29 -2543
rect -29 -3637 29 -3631
rect -29 -3671 -17 -3637
rect -29 -3677 29 -3671
<< nwell >>
rect -211 -3809 211 3809
<< pmos >>
rect -15 2590 15 3590
rect -15 1354 15 2354
rect -15 118 15 1118
rect -15 -1118 15 -118
rect -15 -2354 15 -1354
rect -15 -3590 15 -2590
<< pdiff >>
rect -73 3578 -15 3590
rect -73 2602 -61 3578
rect -27 2602 -15 3578
rect -73 2590 -15 2602
rect 15 3578 73 3590
rect 15 2602 27 3578
rect 61 2602 73 3578
rect 15 2590 73 2602
rect -73 2342 -15 2354
rect -73 1366 -61 2342
rect -27 1366 -15 2342
rect -73 1354 -15 1366
rect 15 2342 73 2354
rect 15 1366 27 2342
rect 61 1366 73 2342
rect 15 1354 73 1366
rect -73 1106 -15 1118
rect -73 130 -61 1106
rect -27 130 -15 1106
rect -73 118 -15 130
rect 15 1106 73 1118
rect 15 130 27 1106
rect 61 130 73 1106
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -1106 -61 -130
rect -27 -1106 -15 -130
rect -73 -1118 -15 -1106
rect 15 -130 73 -118
rect 15 -1106 27 -130
rect 61 -1106 73 -130
rect 15 -1118 73 -1106
rect -73 -1366 -15 -1354
rect -73 -2342 -61 -1366
rect -27 -2342 -15 -1366
rect -73 -2354 -15 -2342
rect 15 -1366 73 -1354
rect 15 -2342 27 -1366
rect 61 -2342 73 -1366
rect 15 -2354 73 -2342
rect -73 -2602 -15 -2590
rect -73 -3578 -61 -2602
rect -27 -3578 -15 -2602
rect -73 -3590 -15 -3578
rect 15 -2602 73 -2590
rect 15 -3578 27 -2602
rect 61 -3578 73 -2602
rect 15 -3590 73 -3578
<< pdiffc >>
rect -61 2602 -27 3578
rect 27 2602 61 3578
rect -61 1366 -27 2342
rect 27 1366 61 2342
rect -61 130 -27 1106
rect 27 130 61 1106
rect -61 -1106 -27 -130
rect 27 -1106 61 -130
rect -61 -2342 -27 -1366
rect 27 -2342 61 -1366
rect -61 -3578 -27 -2602
rect 27 -3578 61 -2602
<< nsubdiff >>
rect -175 3739 -79 3773
rect 79 3739 175 3773
rect -175 3677 -141 3739
rect 141 3677 175 3739
rect -175 -3739 -141 -3677
rect 141 -3739 175 -3677
rect -175 -3773 -79 -3739
rect 79 -3773 175 -3739
<< nsubdiffcont >>
rect -79 3739 79 3773
rect -175 -3677 -141 3677
rect 141 -3677 175 3677
rect -79 -3773 79 -3739
<< poly >>
rect -33 3671 33 3687
rect -33 3637 -17 3671
rect 17 3637 33 3671
rect -33 3621 33 3637
rect -15 3590 15 3621
rect -15 2559 15 2590
rect -33 2543 33 2559
rect -33 2509 -17 2543
rect 17 2509 33 2543
rect -33 2493 33 2509
rect -33 2435 33 2451
rect -33 2401 -17 2435
rect 17 2401 33 2435
rect -33 2385 33 2401
rect -15 2354 15 2385
rect -15 1323 15 1354
rect -33 1307 33 1323
rect -33 1273 -17 1307
rect 17 1273 33 1307
rect -33 1257 33 1273
rect -33 1199 33 1215
rect -33 1165 -17 1199
rect 17 1165 33 1199
rect -33 1149 33 1165
rect -15 1118 15 1149
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -1149 15 -1118
rect -33 -1165 33 -1149
rect -33 -1199 -17 -1165
rect 17 -1199 33 -1165
rect -33 -1215 33 -1199
rect -33 -1273 33 -1257
rect -33 -1307 -17 -1273
rect 17 -1307 33 -1273
rect -33 -1323 33 -1307
rect -15 -1354 15 -1323
rect -15 -2385 15 -2354
rect -33 -2401 33 -2385
rect -33 -2435 -17 -2401
rect 17 -2435 33 -2401
rect -33 -2451 33 -2435
rect -33 -2509 33 -2493
rect -33 -2543 -17 -2509
rect 17 -2543 33 -2509
rect -33 -2559 33 -2543
rect -15 -2590 15 -2559
rect -15 -3621 15 -3590
rect -33 -3637 33 -3621
rect -33 -3671 -17 -3637
rect 17 -3671 33 -3637
rect -33 -3687 33 -3671
<< polycont >>
rect -17 3637 17 3671
rect -17 2509 17 2543
rect -17 2401 17 2435
rect -17 1273 17 1307
rect -17 1165 17 1199
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -1199 17 -1165
rect -17 -1307 17 -1273
rect -17 -2435 17 -2401
rect -17 -2543 17 -2509
rect -17 -3671 17 -3637
<< locali >>
rect -175 3739 -79 3773
rect 79 3739 175 3773
rect -175 3677 -141 3739
rect 141 3677 175 3739
rect -33 3637 -17 3671
rect 17 3637 33 3671
rect -61 3578 -27 3594
rect -61 2586 -27 2602
rect 27 3578 61 3594
rect 27 2586 61 2602
rect -33 2509 -17 2543
rect 17 2509 33 2543
rect -33 2401 -17 2435
rect 17 2401 33 2435
rect -61 2342 -27 2358
rect -61 1350 -27 1366
rect 27 2342 61 2358
rect 27 1350 61 1366
rect -33 1273 -17 1307
rect 17 1273 33 1307
rect -33 1165 -17 1199
rect 17 1165 33 1199
rect -61 1106 -27 1122
rect -61 114 -27 130
rect 27 1106 61 1122
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -1122 -27 -1106
rect 27 -130 61 -114
rect 27 -1122 61 -1106
rect -33 -1199 -17 -1165
rect 17 -1199 33 -1165
rect -33 -1307 -17 -1273
rect 17 -1307 33 -1273
rect -61 -1366 -27 -1350
rect -61 -2358 -27 -2342
rect 27 -1366 61 -1350
rect 27 -2358 61 -2342
rect -33 -2435 -17 -2401
rect 17 -2435 33 -2401
rect -33 -2543 -17 -2509
rect 17 -2543 33 -2509
rect -61 -2602 -27 -2586
rect -61 -3594 -27 -3578
rect 27 -2602 61 -2586
rect 27 -3594 61 -3578
rect -33 -3671 -17 -3637
rect 17 -3671 33 -3637
rect -175 -3739 -141 -3677
rect 141 -3739 175 -3677
rect -175 -3773 -79 -3739
rect 79 -3773 175 -3739
<< viali >>
rect -17 3637 17 3671
rect -61 2602 -27 3578
rect 27 2602 61 3578
rect -17 2509 17 2543
rect -17 2401 17 2435
rect -61 1366 -27 2342
rect 27 1366 61 2342
rect -17 1273 17 1307
rect -17 1165 17 1199
rect -61 130 -27 1106
rect 27 130 61 1106
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -1106 -27 -130
rect 27 -1106 61 -130
rect -17 -1199 17 -1165
rect -17 -1307 17 -1273
rect -61 -2342 -27 -1366
rect 27 -2342 61 -1366
rect -17 -2435 17 -2401
rect -17 -2543 17 -2509
rect -61 -3578 -27 -2602
rect 27 -3578 61 -2602
rect -17 -3671 17 -3637
<< metal1 >>
rect -29 3671 29 3677
rect -29 3637 -17 3671
rect 17 3637 29 3671
rect -29 3631 29 3637
rect -67 3578 -21 3590
rect -67 2602 -61 3578
rect -27 2602 -21 3578
rect -67 2590 -21 2602
rect 21 3578 67 3590
rect 21 2602 27 3578
rect 61 2602 67 3578
rect 21 2590 67 2602
rect -29 2543 29 2549
rect -29 2509 -17 2543
rect 17 2509 29 2543
rect -29 2503 29 2509
rect -29 2435 29 2441
rect -29 2401 -17 2435
rect 17 2401 29 2435
rect -29 2395 29 2401
rect -67 2342 -21 2354
rect -67 1366 -61 2342
rect -27 1366 -21 2342
rect -67 1354 -21 1366
rect 21 2342 67 2354
rect 21 1366 27 2342
rect 61 1366 67 2342
rect 21 1354 67 1366
rect -29 1307 29 1313
rect -29 1273 -17 1307
rect 17 1273 29 1307
rect -29 1267 29 1273
rect -29 1199 29 1205
rect -29 1165 -17 1199
rect 17 1165 29 1199
rect -29 1159 29 1165
rect -67 1106 -21 1118
rect -67 130 -61 1106
rect -27 130 -21 1106
rect -67 118 -21 130
rect 21 1106 67 1118
rect 21 130 27 1106
rect 61 130 67 1106
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -1106 -61 -130
rect -27 -1106 -21 -130
rect -67 -1118 -21 -1106
rect 21 -130 67 -118
rect 21 -1106 27 -130
rect 61 -1106 67 -130
rect 21 -1118 67 -1106
rect -29 -1165 29 -1159
rect -29 -1199 -17 -1165
rect 17 -1199 29 -1165
rect -29 -1205 29 -1199
rect -29 -1273 29 -1267
rect -29 -1307 -17 -1273
rect 17 -1307 29 -1273
rect -29 -1313 29 -1307
rect -67 -1366 -21 -1354
rect -67 -2342 -61 -1366
rect -27 -2342 -21 -1366
rect -67 -2354 -21 -2342
rect 21 -1366 67 -1354
rect 21 -2342 27 -1366
rect 61 -2342 67 -1366
rect 21 -2354 67 -2342
rect -29 -2401 29 -2395
rect -29 -2435 -17 -2401
rect 17 -2435 29 -2401
rect -29 -2441 29 -2435
rect -29 -2509 29 -2503
rect -29 -2543 -17 -2509
rect 17 -2543 29 -2509
rect -29 -2549 29 -2543
rect -67 -2602 -21 -2590
rect -67 -3578 -61 -2602
rect -27 -3578 -21 -2602
rect -67 -3590 -21 -3578
rect 21 -2602 67 -2590
rect 21 -3578 27 -2602
rect 61 -3578 67 -2602
rect 21 -3590 67 -3578
rect -29 -3637 29 -3631
rect -29 -3671 -17 -3637
rect 17 -3671 29 -3637
rect -29 -3677 29 -3671
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -158 -3756 158 3756
string parameters w 5 l 0.15 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
