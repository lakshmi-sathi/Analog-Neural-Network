magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_s >>
rect 14540 -1351 14898 -1282
rect 14708 -1450 14730 -1351
rect 14804 -1450 14898 -1351
rect 14708 -1451 14898 -1450
rect 14672 -1557 14898 -1451
rect 14672 -1595 14766 -1557
rect 14804 -1595 14898 -1557
rect 14672 -1619 14898 -1595
rect 14548 -2605 14906 -2536
rect 14716 -2704 14738 -2605
rect 14812 -2704 14906 -2605
rect 14716 -2705 14906 -2704
rect 14680 -2811 14906 -2705
rect 14680 -2849 14774 -2811
rect 14812 -2849 14906 -2811
rect 14680 -2873 14906 -2849
rect 14528 -3873 14886 -3804
rect 14696 -3972 14718 -3873
rect 14792 -3972 14886 -3873
rect 14696 -3973 14886 -3972
rect 14660 -4079 14886 -3973
rect 14660 -4117 14754 -4079
rect 14792 -4117 14886 -4079
rect 14660 -4141 14886 -4117
<< locali >>
rect 14006 -1292 14420 -1200
rect 14014 -2542 14428 -2450
rect 13992 -3810 14406 -3718
<< metal1 >>
rect 586 2556 1016 2578
rect 582 2532 1016 2556
rect 582 2096 607 2532
rect 979 2096 1016 2532
rect 582 2072 1016 2096
rect 586 1944 1016 2072
rect -514 1402 1016 1944
rect 586 1184 1016 1402
rect 11922 1672 12160 1674
rect 11922 1086 12374 1672
rect 12114 -1102 12374 1086
rect 13838 1550 15688 1910
rect 13838 -328 14198 1550
rect 15328 1208 15688 1550
rect 26632 1201 27262 1208
rect 26632 957 26667 1201
rect 27231 957 27262 1201
rect 26632 950 27262 957
rect 13838 -688 18768 -328
rect 614 -1498 956 -1222
rect -540 -2040 956 -1498
rect 11890 -1692 12374 -1102
rect 614 -2226 956 -2040
rect 614 -2254 966 -2226
rect 614 -2562 637 -2254
rect 945 -2562 966 -2254
rect 614 -2590 966 -2562
rect 614 -2604 956 -2590
rect 12114 -2942 12374 -1692
rect 14834 -1584 15196 -1565
rect 18370 -1566 18730 -688
rect 14834 -1764 14845 -1584
rect 14961 -1764 15196 -1584
rect 14834 -1787 15196 -1764
rect 18270 -1788 18730 -1566
rect 18298 -1790 18730 -1788
rect 18370 -2768 18730 -1790
rect 14840 -2818 15210 -2810
rect 14836 -2825 15210 -2818
rect 12114 -2964 13044 -2942
rect 12114 -3656 12498 -2964
rect 12998 -3108 13044 -2964
rect 14836 -3005 14851 -2825
rect 14967 -3005 15210 -2825
rect 18270 -2990 18730 -2768
rect 14836 -3012 15210 -3005
rect 14840 -3022 15210 -3012
rect 12998 -3336 13040 -3108
rect 12998 -3656 13044 -3336
rect 12114 -3668 13044 -3656
rect 600 -3857 926 -3830
rect 600 -4165 643 -3857
rect 887 -4165 926 -3857
rect 600 -4306 926 -4165
rect -548 -4848 936 -4306
rect 12114 -4584 12374 -3668
rect 18370 -4048 18730 -2990
rect 20194 -2776 20552 -2768
rect 20194 -3852 20219 -2776
rect 20527 -3852 20552 -2776
rect 20194 -3888 20552 -3852
rect 14828 -4084 15202 -4078
rect 14818 -4092 15202 -4084
rect 14818 -4272 14830 -4092
rect 14946 -4272 15202 -4092
rect 18272 -4266 18730 -4048
rect 14818 -4280 15202 -4272
rect 18370 -4284 18730 -4266
rect 600 -5180 926 -4848
rect 11944 -5132 12374 -4584
rect 12114 -5136 12374 -5132
<< via1 >>
rect 607 2096 979 2532
rect 26667 957 27231 1201
rect 637 -2562 945 -2254
rect 14845 -1764 14961 -1584
rect 12498 -3656 12998 -2964
rect 14851 -3005 14967 -2825
rect 643 -4165 887 -3857
rect 20219 -3852 20527 -2776
rect 14830 -4272 14946 -4092
<< metal2 >>
rect 376 3148 29806 3151
rect 92 3021 30028 3148
rect 92 3014 1595 3021
rect 94 -2996 350 3014
rect 26040 2967 30028 3021
rect 592 2542 994 2566
rect 592 2086 605 2542
rect 981 2086 994 2542
rect 592 2062 994 2086
rect 26652 1201 27246 1212
rect 26652 957 26667 1201
rect 27231 1187 27246 1201
rect 27242 971 27246 1187
rect 27231 957 27246 971
rect 26652 946 27246 957
rect 1399 28 26795 130
rect 1399 -108 19056 28
rect 21112 -108 26795 28
rect 1399 -112 26795 -108
rect 19024 -138 21144 -112
rect 19312 -414 20022 -412
rect 29622 -414 30028 2967
rect 19312 -590 30028 -414
rect 14718 -734 30028 -590
rect 14718 -777 20022 -734
rect 14708 -859 20022 -777
rect 14708 -1402 14790 -859
rect 14828 -1584 14974 -1559
rect 14828 -1764 14845 -1584
rect 14961 -1764 14974 -1584
rect 14828 -1789 14974 -1764
rect 626 -2254 956 -2216
rect 626 -2562 637 -2254
rect 945 -2562 956 -2254
rect 17121 -2313 17203 -859
rect 626 -2600 956 -2562
rect 14711 -2395 17203 -2313
rect 14711 -2649 14793 -2395
rect 14846 -2810 14972 -2808
rect 14838 -2825 14984 -2810
rect 12460 -2964 13056 -2940
rect 94 -3252 11994 -2996
rect 12460 -3108 12498 -2964
rect 12462 -3336 12498 -3108
rect 12460 -3656 12498 -3336
rect 12998 -3656 13056 -2964
rect 14838 -3005 14851 -2825
rect 14967 -3005 14984 -2825
rect 14838 -3020 14984 -3005
rect 14846 -3022 14972 -3020
rect 18659 -3507 18741 -859
rect 19312 -866 20022 -859
rect 20212 -2776 20534 -2758
rect 20212 -2940 20219 -2776
rect 12460 -3670 13056 -3656
rect 616 -3857 914 -3826
rect 616 -3863 643 -3857
rect 887 -3863 914 -3857
rect 616 -4159 617 -3863
rect 913 -4159 914 -3863
rect 12473 -4032 13056 -3670
rect 14689 -3589 18741 -3507
rect 14689 -3925 14771 -3589
rect 19212 -3670 20219 -2940
rect 616 -4165 643 -4159
rect 887 -4165 914 -4159
rect 616 -4196 914 -4165
rect 12472 -4304 13056 -4032
rect 14828 -4080 14948 -4074
rect 14820 -4092 14958 -4080
rect 14820 -4272 14830 -4092
rect 14946 -4272 14958 -4092
rect 14820 -4284 14958 -4272
rect 14828 -4290 14948 -4284
rect 12473 -4900 13056 -4304
rect 12473 -5148 13048 -4900
rect 19212 -5148 19815 -3670
rect 20212 -3852 20219 -3670
rect 20527 -2940 20534 -2776
rect 20527 -2958 27437 -2940
rect 20527 -3654 26723 -2958
rect 27419 -3654 27437 -2958
rect 20527 -3670 27437 -3654
rect 20527 -3852 20534 -3670
rect 20212 -3870 20534 -3852
rect 12473 -5697 19815 -5148
rect 19218 -6000 19910 -5966
rect 27612 -6000 28408 -5822
rect 19212 -6092 19256 -6000
rect 1616 -6216 19256 -6092
rect 19872 -6092 28408 -6000
rect 19872 -6216 28431 -6092
rect 1616 -6266 28431 -6216
<< via2 >>
rect 605 2532 981 2542
rect 605 2096 607 2532
rect 607 2096 979 2532
rect 979 2096 981 2532
rect 605 2086 981 2096
rect 26946 971 27231 1187
rect 27231 971 27242 1187
rect 19056 -108 21112 28
rect 643 -2556 939 -2260
rect 617 -4159 643 -3863
rect 643 -4159 887 -3863
rect 887 -4159 913 -3863
rect 20225 -3822 20521 -2806
rect 26723 -3654 27419 -2958
rect 19256 -6216 19872 -6000
<< metal3 >>
rect 582 2546 1004 2561
rect 582 2082 601 2546
rect 985 2082 1004 2546
rect 582 2067 1004 2082
rect 26920 1187 27276 1214
rect 26920 971 26946 1187
rect 27242 971 27276 1187
rect 11868 166 13582 486
rect 11862 -474 12740 -154
rect 616 -2256 966 -2221
rect 616 -2560 639 -2256
rect 943 -2560 966 -2256
rect 616 -2595 966 -2560
rect 12420 -3008 12740 -474
rect 13262 -1468 13582 166
rect 19000 28 21164 56
rect 19000 -108 19056 28
rect 21112 -108 21164 28
rect 19000 -136 21164 -108
rect 13262 -1750 13578 -1468
rect 13262 -1756 13670 -1750
rect 13262 -1757 13774 -1756
rect 13262 -1854 13944 -1757
rect 13774 -1855 13944 -1854
rect 13614 -3008 13962 -3006
rect 12420 -3108 13962 -3008
rect 606 -3859 924 -3831
rect 606 -3863 653 -3859
rect 877 -3863 924 -3859
rect 606 -4159 617 -3863
rect 913 -4159 924 -3863
rect 606 -4163 653 -4159
rect 877 -4163 924 -4159
rect 606 -4191 924 -4163
rect 12440 -4274 12760 -4272
rect 13776 -4274 13938 -4273
rect 12440 -4367 13938 -4274
rect 12440 -4368 13780 -4367
rect 12440 -5764 12760 -4368
rect 11882 -6084 12760 -5764
rect 19218 -5971 19914 -136
rect 20202 -2806 20544 -2763
rect 20202 -3822 20225 -2806
rect 20521 -3822 20544 -2806
rect 26920 -2949 27276 971
rect 26712 -2958 27430 -2949
rect 26712 -3654 26723 -2958
rect 27419 -3654 27430 -2958
rect 26712 -3663 27430 -3654
rect 20202 -3865 20544 -3822
rect 19208 -6000 19920 -5971
rect 19208 -6216 19256 -6000
rect 19872 -6216 19920 -6000
rect 19208 -6245 19920 -6216
<< via3 >>
rect 601 2542 985 2546
rect 601 2086 605 2542
rect 605 2086 981 2542
rect 981 2086 985 2542
rect 601 2082 985 2086
rect 639 -2260 943 -2256
rect 639 -2556 643 -2260
rect 643 -2556 939 -2260
rect 939 -2556 943 -2260
rect 639 -2560 943 -2556
rect 653 -3863 877 -3859
rect 653 -4159 877 -3863
rect 653 -4163 877 -4159
<< metal4 >>
rect 574 2546 13176 2580
rect 574 2082 601 2546
rect 985 2196 13176 2546
rect 985 2082 1016 2196
rect 574 2054 1016 2082
rect 12792 -1472 13176 2196
rect 30232 1966 30658 2134
rect 30188 1960 30658 1966
rect 27450 1505 30658 1960
rect 27450 1185 28143 1505
rect 30188 1504 30658 1505
rect 30232 1372 30658 1504
rect 12792 -1592 13956 -1472
rect 13278 -2224 13406 -2222
rect 610 -2256 13406 -2224
rect 610 -2560 639 -2256
rect 943 -2560 13406 -2256
rect 610 -2608 13406 -2560
rect 12938 -2614 13406 -2608
rect 13100 -2704 13406 -2614
rect 13100 -2832 13960 -2704
rect 13100 -2834 13352 -2832
rect 582 -3859 12916 -3818
rect 582 -4163 653 -3859
rect 877 -4006 12916 -3859
rect 877 -4104 13934 -4006
rect 877 -4163 12916 -4104
rect 582 -4202 12916 -4163
use mux  mux_2
timestamp 1627926120
transform 1 0 13834 0 -1 -4119
box -22 -348 1124 429
use mux  mux_1
timestamp 1627926120
transform 1 0 13854 0 -1 -2851
box -22 -348 1124 429
use mux  mux_0
timestamp 1627926120
transform 1 0 13846 0 -1 -1597
box -22 -348 1124 429
use voltage_div  voltage_div_0
timestamp 1627926120
transform 1 0 20412 0 1 -3066
box 0 -2992 8012 2542
use analogneuron_invopamp_re_15kfeedbck  analogneuron_invopamp_re_15kfeedbck_0
timestamp 1627926120
transform 1 0 1354 0 1 234
box -1354 -234 10724 2910
use analogneuron_invopamp_re_15kfeedbck  analogneuron_invopamp_re_15kfeedbck_1
timestamp 1627926120
transform 1 0 1348 0 -1 -216
box -1354 -234 10724 2910
use analogneuron_invopamp_re_15kfeedbck  analogneuron_invopamp_re_15kfeedbck_2
timestamp 1627926120
transform 1 0 1358 0 1 -6032
box -1354 -234 10724 2910
use analogneuron_invopamp_re_15kfeedbck_ReLU  analogneuron_invopamp_re_15kfeedbck_ReLU_0
timestamp 1627926120
transform 1 0 16082 0 1 241
box -1354 -343 13246 2910
<< labels >>
rlabel metal1 s 15048 -1772 15184 -1574 4 r1p1
port 1 nsew
rlabel metal1 s 15068 -3012 15204 -2814 4 r2p1
port 2 nsew
rlabel metal1 s 15052 -4278 15188 -4080 4 r3p1
port 3 nsew
rlabel metal1 s 18288 -4256 18424 -4058 4 r3p2
port 4 nsew
rlabel metal2 s 1366 3026 30014 3140 4 VDD
port 5 nsew
rlabel metal2 s 1444 -3244 11944 -3020 4 VDD
port 5 nsew
rlabel metal2 s 1626 -6256 28406 -6126 4 GND
port 6 nsew
rlabel metal2 s 1414 -90 12030 118 4 GND
port 6 nsew
rlabel locali s 13998 -3804 14394 -3730 4 m3sel
port 7 nsew
rlabel locali s 14022 -2534 14418 -2460 4 m2sel
port 8 nsew
rlabel locali s 14012 -1282 14408 -1208 4 m1sel
port 9 nsew
rlabel metal1 s -492 1428 -86 1922 4 in1
port 10 nsew
rlabel metal1 s -514 -2020 -108 -1526 4 in2
port 11 nsew
rlabel metal1 s -516 -4822 -110 -4328 4 in3
port 12 nsew
rlabel metal4 s 30250 1384 30628 2108 4 out
port 13 nsew
rlabel metal2 s 12482 -3690 13028 -2954 4 vcm
port 14 nsew
<< end >>
