magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 99 35 531
rect -35 -531 35 -99
<< xpolyres >>
rect -35 -99 35 99
<< viali >>
rect -17 477 17 511
rect -17 405 17 439
rect -17 333 17 367
rect -17 261 17 295
rect -17 189 17 223
rect -17 117 17 151
rect -17 -152 17 -118
rect -17 -224 17 -190
rect -17 -296 17 -262
rect -17 -368 17 -334
rect -17 -440 17 -406
rect -17 -512 17 -478
<< metal1 >>
rect -25 511 25 525
rect -25 477 -17 511
rect 17 477 25 511
rect -25 439 25 477
rect -25 405 -17 439
rect 17 405 25 439
rect -25 367 25 405
rect -25 333 -17 367
rect 17 333 25 367
rect -25 295 25 333
rect -25 261 -17 295
rect 17 261 25 295
rect -25 223 25 261
rect -25 189 -17 223
rect 17 189 25 223
rect -25 151 25 189
rect -25 117 -17 151
rect 17 117 25 151
rect -25 104 25 117
rect -25 -118 25 -104
rect -25 -152 -17 -118
rect 17 -152 25 -118
rect -25 -190 25 -152
rect -25 -224 -17 -190
rect 17 -224 25 -190
rect -25 -262 25 -224
rect -25 -296 -17 -262
rect 17 -296 25 -262
rect -25 -334 25 -296
rect -25 -368 -17 -334
rect 17 -368 25 -334
rect -25 -406 25 -368
rect -25 -440 -17 -406
rect 17 -440 25 -406
rect -25 -478 25 -440
rect -25 -512 -17 -478
rect 17 -512 25 -478
rect -25 -525 25 -512
<< end >>
