magic
tech sky130A
magscale 1 2
timestamp 1628375762
<< xpolycontact >>
rect -69 210 69 642
rect -69 -642 69 -210
<< ppolyres >>
rect -69 -210 69 210
<< viali >>
rect -53 227 53 624
rect -53 -624 53 -227
<< metal1 >>
rect -59 624 59 636
rect -59 227 -53 624
rect 53 227 59 624
rect -59 215 59 227
rect -59 -227 59 -215
rect -59 -624 -53 -227
rect 53 -624 59 -227
rect -59 -636 59 -624
<< res0p69 >>
rect -71 -212 71 212
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p69
string parameters w 0.690 l 2.1 m 1 nx 1 wmin 0.690 lmin 0.50 rho 319.8 val 1.028k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
