magic
tech sky130A
magscale 1 2
timestamp 1627923075
<< xpolycontact >>
rect -35 605 35 1037
rect -35 -1037 35 -605
<< ppolyres >>
rect -35 -605 35 605
<< viali >>
rect -19 622 19 1019
rect -19 -1019 19 -622
<< metal1 >>
rect -25 1019 25 1031
rect -25 622 -19 1019
rect 19 622 25 1019
rect -25 610 25 622
rect -25 -622 25 -610
rect -25 -1019 -19 -622
rect 19 -1019 25 -622
rect -25 -1031 25 -1019
<< res0p35 >>
rect -37 -607 37 607
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string parameters w 0.350 l 6.05 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 5.637k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 0.350 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
