magic
tech sky130A
magscale 1 2
timestamp 1626800441
<< error_p >>
rect -1901 372 -1843 378
rect -1709 372 -1651 378
rect -1517 372 -1459 378
rect -1325 372 -1267 378
rect -1133 372 -1075 378
rect -941 372 -883 378
rect -749 372 -691 378
rect -557 372 -499 378
rect -365 372 -307 378
rect -173 372 -115 378
rect 19 372 77 378
rect 211 372 269 378
rect 403 372 461 378
rect 595 372 653 378
rect 787 372 845 378
rect 979 372 1037 378
rect 1171 372 1229 378
rect 1363 372 1421 378
rect 1555 372 1613 378
rect 1747 372 1805 378
rect 1939 372 1997 378
rect -1901 338 -1889 372
rect -1709 338 -1697 372
rect -1517 338 -1505 372
rect -1325 338 -1313 372
rect -1133 338 -1121 372
rect -941 338 -929 372
rect -749 338 -737 372
rect -557 338 -545 372
rect -365 338 -353 372
rect -173 338 -161 372
rect 19 338 31 372
rect 211 338 223 372
rect 403 338 415 372
rect 595 338 607 372
rect 787 338 799 372
rect 979 338 991 372
rect 1171 338 1183 372
rect 1363 338 1375 372
rect 1555 338 1567 372
rect 1747 338 1759 372
rect 1939 338 1951 372
rect -1901 332 -1843 338
rect -1709 332 -1651 338
rect -1517 332 -1459 338
rect -1325 332 -1267 338
rect -1133 332 -1075 338
rect -941 332 -883 338
rect -749 332 -691 338
rect -557 332 -499 338
rect -365 332 -307 338
rect -173 332 -115 338
rect 19 332 77 338
rect 211 332 269 338
rect 403 332 461 338
rect 595 332 653 338
rect 787 332 845 338
rect 979 332 1037 338
rect 1171 332 1229 338
rect 1363 332 1421 338
rect 1555 332 1613 338
rect 1747 332 1805 338
rect 1939 332 1997 338
rect -1997 -338 -1939 -332
rect -1805 -338 -1747 -332
rect -1613 -338 -1555 -332
rect -1421 -338 -1363 -332
rect -1229 -338 -1171 -332
rect -1037 -338 -979 -332
rect -845 -338 -787 -332
rect -653 -338 -595 -332
rect -461 -338 -403 -332
rect -269 -338 -211 -332
rect -77 -338 -19 -332
rect 115 -338 173 -332
rect 307 -338 365 -332
rect 499 -338 557 -332
rect 691 -338 749 -332
rect 883 -338 941 -332
rect 1075 -338 1133 -332
rect 1267 -338 1325 -332
rect 1459 -338 1517 -332
rect 1651 -338 1709 -332
rect 1843 -338 1901 -332
rect -1997 -372 -1985 -338
rect -1805 -372 -1793 -338
rect -1613 -372 -1601 -338
rect -1421 -372 -1409 -338
rect -1229 -372 -1217 -338
rect -1037 -372 -1025 -338
rect -845 -372 -833 -338
rect -653 -372 -641 -338
rect -461 -372 -449 -338
rect -269 -372 -257 -338
rect -77 -372 -65 -338
rect 115 -372 127 -338
rect 307 -372 319 -338
rect 499 -372 511 -338
rect 691 -372 703 -338
rect 883 -372 895 -338
rect 1075 -372 1087 -338
rect 1267 -372 1279 -338
rect 1459 -372 1471 -338
rect 1651 -372 1663 -338
rect 1843 -372 1855 -338
rect -1997 -378 -1939 -372
rect -1805 -378 -1747 -372
rect -1613 -378 -1555 -372
rect -1421 -378 -1363 -372
rect -1229 -378 -1171 -372
rect -1037 -378 -979 -372
rect -845 -378 -787 -372
rect -653 -378 -595 -372
rect -461 -378 -403 -372
rect -269 -378 -211 -372
rect -77 -378 -19 -372
rect 115 -378 173 -372
rect 307 -378 365 -372
rect 499 -378 557 -372
rect 691 -378 749 -372
rect 883 -378 941 -372
rect 1075 -378 1133 -372
rect 1267 -378 1325 -372
rect 1459 -378 1517 -372
rect 1651 -378 1709 -372
rect 1843 -378 1901 -372
<< pwell >>
rect -2183 -510 2183 510
<< nmos >>
rect -1983 -300 -1953 300
rect -1887 -300 -1857 300
rect -1791 -300 -1761 300
rect -1695 -300 -1665 300
rect -1599 -300 -1569 300
rect -1503 -300 -1473 300
rect -1407 -300 -1377 300
rect -1311 -300 -1281 300
rect -1215 -300 -1185 300
rect -1119 -300 -1089 300
rect -1023 -300 -993 300
rect -927 -300 -897 300
rect -831 -300 -801 300
rect -735 -300 -705 300
rect -639 -300 -609 300
rect -543 -300 -513 300
rect -447 -300 -417 300
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
rect 417 -300 447 300
rect 513 -300 543 300
rect 609 -300 639 300
rect 705 -300 735 300
rect 801 -300 831 300
rect 897 -300 927 300
rect 993 -300 1023 300
rect 1089 -300 1119 300
rect 1185 -300 1215 300
rect 1281 -300 1311 300
rect 1377 -300 1407 300
rect 1473 -300 1503 300
rect 1569 -300 1599 300
rect 1665 -300 1695 300
rect 1761 -300 1791 300
rect 1857 -300 1887 300
rect 1953 -300 1983 300
<< ndiff >>
rect -2045 288 -1983 300
rect -2045 -288 -2033 288
rect -1999 -288 -1983 288
rect -2045 -300 -1983 -288
rect -1953 288 -1887 300
rect -1953 -288 -1937 288
rect -1903 -288 -1887 288
rect -1953 -300 -1887 -288
rect -1857 288 -1791 300
rect -1857 -288 -1841 288
rect -1807 -288 -1791 288
rect -1857 -300 -1791 -288
rect -1761 288 -1695 300
rect -1761 -288 -1745 288
rect -1711 -288 -1695 288
rect -1761 -300 -1695 -288
rect -1665 288 -1599 300
rect -1665 -288 -1649 288
rect -1615 -288 -1599 288
rect -1665 -300 -1599 -288
rect -1569 288 -1503 300
rect -1569 -288 -1553 288
rect -1519 -288 -1503 288
rect -1569 -300 -1503 -288
rect -1473 288 -1407 300
rect -1473 -288 -1457 288
rect -1423 -288 -1407 288
rect -1473 -300 -1407 -288
rect -1377 288 -1311 300
rect -1377 -288 -1361 288
rect -1327 -288 -1311 288
rect -1377 -300 -1311 -288
rect -1281 288 -1215 300
rect -1281 -288 -1265 288
rect -1231 -288 -1215 288
rect -1281 -300 -1215 -288
rect -1185 288 -1119 300
rect -1185 -288 -1169 288
rect -1135 -288 -1119 288
rect -1185 -300 -1119 -288
rect -1089 288 -1023 300
rect -1089 -288 -1073 288
rect -1039 -288 -1023 288
rect -1089 -300 -1023 -288
rect -993 288 -927 300
rect -993 -288 -977 288
rect -943 -288 -927 288
rect -993 -300 -927 -288
rect -897 288 -831 300
rect -897 -288 -881 288
rect -847 -288 -831 288
rect -897 -300 -831 -288
rect -801 288 -735 300
rect -801 -288 -785 288
rect -751 -288 -735 288
rect -801 -300 -735 -288
rect -705 288 -639 300
rect -705 -288 -689 288
rect -655 -288 -639 288
rect -705 -300 -639 -288
rect -609 288 -543 300
rect -609 -288 -593 288
rect -559 -288 -543 288
rect -609 -300 -543 -288
rect -513 288 -447 300
rect -513 -288 -497 288
rect -463 -288 -447 288
rect -513 -300 -447 -288
rect -417 288 -351 300
rect -417 -288 -401 288
rect -367 -288 -351 288
rect -417 -300 -351 -288
rect -321 288 -255 300
rect -321 -288 -305 288
rect -271 -288 -255 288
rect -321 -300 -255 -288
rect -225 288 -159 300
rect -225 -288 -209 288
rect -175 -288 -159 288
rect -225 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 225 300
rect 159 -288 175 288
rect 209 -288 225 288
rect 159 -300 225 -288
rect 255 288 321 300
rect 255 -288 271 288
rect 305 -288 321 288
rect 255 -300 321 -288
rect 351 288 417 300
rect 351 -288 367 288
rect 401 -288 417 288
rect 351 -300 417 -288
rect 447 288 513 300
rect 447 -288 463 288
rect 497 -288 513 288
rect 447 -300 513 -288
rect 543 288 609 300
rect 543 -288 559 288
rect 593 -288 609 288
rect 543 -300 609 -288
rect 639 288 705 300
rect 639 -288 655 288
rect 689 -288 705 288
rect 639 -300 705 -288
rect 735 288 801 300
rect 735 -288 751 288
rect 785 -288 801 288
rect 735 -300 801 -288
rect 831 288 897 300
rect 831 -288 847 288
rect 881 -288 897 288
rect 831 -300 897 -288
rect 927 288 993 300
rect 927 -288 943 288
rect 977 -288 993 288
rect 927 -300 993 -288
rect 1023 288 1089 300
rect 1023 -288 1039 288
rect 1073 -288 1089 288
rect 1023 -300 1089 -288
rect 1119 288 1185 300
rect 1119 -288 1135 288
rect 1169 -288 1185 288
rect 1119 -300 1185 -288
rect 1215 288 1281 300
rect 1215 -288 1231 288
rect 1265 -288 1281 288
rect 1215 -300 1281 -288
rect 1311 288 1377 300
rect 1311 -288 1327 288
rect 1361 -288 1377 288
rect 1311 -300 1377 -288
rect 1407 288 1473 300
rect 1407 -288 1423 288
rect 1457 -288 1473 288
rect 1407 -300 1473 -288
rect 1503 288 1569 300
rect 1503 -288 1519 288
rect 1553 -288 1569 288
rect 1503 -300 1569 -288
rect 1599 288 1665 300
rect 1599 -288 1615 288
rect 1649 -288 1665 288
rect 1599 -300 1665 -288
rect 1695 288 1761 300
rect 1695 -288 1711 288
rect 1745 -288 1761 288
rect 1695 -300 1761 -288
rect 1791 288 1857 300
rect 1791 -288 1807 288
rect 1841 -288 1857 288
rect 1791 -300 1857 -288
rect 1887 288 1953 300
rect 1887 -288 1903 288
rect 1937 -288 1953 288
rect 1887 -300 1953 -288
rect 1983 288 2045 300
rect 1983 -288 1999 288
rect 2033 -288 2045 288
rect 1983 -300 2045 -288
<< ndiffc >>
rect -2033 -288 -1999 288
rect -1937 -288 -1903 288
rect -1841 -288 -1807 288
rect -1745 -288 -1711 288
rect -1649 -288 -1615 288
rect -1553 -288 -1519 288
rect -1457 -288 -1423 288
rect -1361 -288 -1327 288
rect -1265 -288 -1231 288
rect -1169 -288 -1135 288
rect -1073 -288 -1039 288
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
rect 1039 -288 1073 288
rect 1135 -288 1169 288
rect 1231 -288 1265 288
rect 1327 -288 1361 288
rect 1423 -288 1457 288
rect 1519 -288 1553 288
rect 1615 -288 1649 288
rect 1711 -288 1745 288
rect 1807 -288 1841 288
rect 1903 -288 1937 288
rect 1999 -288 2033 288
<< psubdiff >>
rect -2147 440 -2051 474
rect 2051 440 2147 474
rect -2147 378 -2113 440
rect 2113 378 2147 440
rect -2147 -440 -2113 -378
rect 2113 -440 2147 -378
rect -2147 -474 -2051 -440
rect 2051 -474 2147 -440
<< psubdiffcont >>
rect -2051 440 2051 474
rect -2147 -378 -2113 378
rect 2113 -378 2147 378
rect -2051 -474 2051 -440
<< poly >>
rect -1905 372 -1839 388
rect -1905 338 -1889 372
rect -1855 338 -1839 372
rect -1983 300 -1953 326
rect -1905 322 -1839 338
rect -1713 372 -1647 388
rect -1713 338 -1697 372
rect -1663 338 -1647 372
rect -1887 300 -1857 322
rect -1791 300 -1761 326
rect -1713 322 -1647 338
rect -1521 372 -1455 388
rect -1521 338 -1505 372
rect -1471 338 -1455 372
rect -1695 300 -1665 322
rect -1599 300 -1569 326
rect -1521 322 -1455 338
rect -1329 372 -1263 388
rect -1329 338 -1313 372
rect -1279 338 -1263 372
rect -1503 300 -1473 322
rect -1407 300 -1377 326
rect -1329 322 -1263 338
rect -1137 372 -1071 388
rect -1137 338 -1121 372
rect -1087 338 -1071 372
rect -1311 300 -1281 322
rect -1215 300 -1185 326
rect -1137 322 -1071 338
rect -945 372 -879 388
rect -945 338 -929 372
rect -895 338 -879 372
rect -1119 300 -1089 322
rect -1023 300 -993 326
rect -945 322 -879 338
rect -753 372 -687 388
rect -753 338 -737 372
rect -703 338 -687 372
rect -927 300 -897 322
rect -831 300 -801 326
rect -753 322 -687 338
rect -561 372 -495 388
rect -561 338 -545 372
rect -511 338 -495 372
rect -735 300 -705 322
rect -639 300 -609 326
rect -561 322 -495 338
rect -369 372 -303 388
rect -369 338 -353 372
rect -319 338 -303 372
rect -543 300 -513 322
rect -447 300 -417 326
rect -369 322 -303 338
rect -177 372 -111 388
rect -177 338 -161 372
rect -127 338 -111 372
rect -351 300 -321 322
rect -255 300 -225 326
rect -177 322 -111 338
rect 15 372 81 388
rect 15 338 31 372
rect 65 338 81 372
rect -159 300 -129 322
rect -63 300 -33 326
rect 15 322 81 338
rect 207 372 273 388
rect 207 338 223 372
rect 257 338 273 372
rect 33 300 63 322
rect 129 300 159 326
rect 207 322 273 338
rect 399 372 465 388
rect 399 338 415 372
rect 449 338 465 372
rect 225 300 255 322
rect 321 300 351 326
rect 399 322 465 338
rect 591 372 657 388
rect 591 338 607 372
rect 641 338 657 372
rect 417 300 447 322
rect 513 300 543 326
rect 591 322 657 338
rect 783 372 849 388
rect 783 338 799 372
rect 833 338 849 372
rect 609 300 639 322
rect 705 300 735 326
rect 783 322 849 338
rect 975 372 1041 388
rect 975 338 991 372
rect 1025 338 1041 372
rect 801 300 831 322
rect 897 300 927 326
rect 975 322 1041 338
rect 1167 372 1233 388
rect 1167 338 1183 372
rect 1217 338 1233 372
rect 993 300 1023 322
rect 1089 300 1119 326
rect 1167 322 1233 338
rect 1359 372 1425 388
rect 1359 338 1375 372
rect 1409 338 1425 372
rect 1185 300 1215 322
rect 1281 300 1311 326
rect 1359 322 1425 338
rect 1551 372 1617 388
rect 1551 338 1567 372
rect 1601 338 1617 372
rect 1377 300 1407 322
rect 1473 300 1503 326
rect 1551 322 1617 338
rect 1743 372 1809 388
rect 1743 338 1759 372
rect 1793 338 1809 372
rect 1569 300 1599 322
rect 1665 300 1695 326
rect 1743 322 1809 338
rect 1935 372 2001 388
rect 1935 338 1951 372
rect 1985 338 2001 372
rect 1761 300 1791 322
rect 1857 300 1887 326
rect 1935 322 2001 338
rect 1953 300 1983 322
rect -1983 -322 -1953 -300
rect -2001 -338 -1935 -322
rect -1887 -326 -1857 -300
rect -1791 -322 -1761 -300
rect -2001 -372 -1985 -338
rect -1951 -372 -1935 -338
rect -2001 -388 -1935 -372
rect -1809 -338 -1743 -322
rect -1695 -326 -1665 -300
rect -1599 -322 -1569 -300
rect -1809 -372 -1793 -338
rect -1759 -372 -1743 -338
rect -1809 -388 -1743 -372
rect -1617 -338 -1551 -322
rect -1503 -326 -1473 -300
rect -1407 -322 -1377 -300
rect -1617 -372 -1601 -338
rect -1567 -372 -1551 -338
rect -1617 -388 -1551 -372
rect -1425 -338 -1359 -322
rect -1311 -326 -1281 -300
rect -1215 -322 -1185 -300
rect -1425 -372 -1409 -338
rect -1375 -372 -1359 -338
rect -1425 -388 -1359 -372
rect -1233 -338 -1167 -322
rect -1119 -326 -1089 -300
rect -1023 -322 -993 -300
rect -1233 -372 -1217 -338
rect -1183 -372 -1167 -338
rect -1233 -388 -1167 -372
rect -1041 -338 -975 -322
rect -927 -326 -897 -300
rect -831 -322 -801 -300
rect -1041 -372 -1025 -338
rect -991 -372 -975 -338
rect -1041 -388 -975 -372
rect -849 -338 -783 -322
rect -735 -326 -705 -300
rect -639 -322 -609 -300
rect -849 -372 -833 -338
rect -799 -372 -783 -338
rect -849 -388 -783 -372
rect -657 -338 -591 -322
rect -543 -326 -513 -300
rect -447 -322 -417 -300
rect -657 -372 -641 -338
rect -607 -372 -591 -338
rect -657 -388 -591 -372
rect -465 -338 -399 -322
rect -351 -326 -321 -300
rect -255 -322 -225 -300
rect -465 -372 -449 -338
rect -415 -372 -399 -338
rect -465 -388 -399 -372
rect -273 -338 -207 -322
rect -159 -326 -129 -300
rect -63 -322 -33 -300
rect -273 -372 -257 -338
rect -223 -372 -207 -338
rect -273 -388 -207 -372
rect -81 -338 -15 -322
rect 33 -326 63 -300
rect 129 -322 159 -300
rect -81 -372 -65 -338
rect -31 -372 -15 -338
rect -81 -388 -15 -372
rect 111 -338 177 -322
rect 225 -326 255 -300
rect 321 -322 351 -300
rect 111 -372 127 -338
rect 161 -372 177 -338
rect 111 -388 177 -372
rect 303 -338 369 -322
rect 417 -326 447 -300
rect 513 -322 543 -300
rect 303 -372 319 -338
rect 353 -372 369 -338
rect 303 -388 369 -372
rect 495 -338 561 -322
rect 609 -326 639 -300
rect 705 -322 735 -300
rect 495 -372 511 -338
rect 545 -372 561 -338
rect 495 -388 561 -372
rect 687 -338 753 -322
rect 801 -326 831 -300
rect 897 -322 927 -300
rect 687 -372 703 -338
rect 737 -372 753 -338
rect 687 -388 753 -372
rect 879 -338 945 -322
rect 993 -326 1023 -300
rect 1089 -322 1119 -300
rect 879 -372 895 -338
rect 929 -372 945 -338
rect 879 -388 945 -372
rect 1071 -338 1137 -322
rect 1185 -326 1215 -300
rect 1281 -322 1311 -300
rect 1071 -372 1087 -338
rect 1121 -372 1137 -338
rect 1071 -388 1137 -372
rect 1263 -338 1329 -322
rect 1377 -326 1407 -300
rect 1473 -322 1503 -300
rect 1263 -372 1279 -338
rect 1313 -372 1329 -338
rect 1263 -388 1329 -372
rect 1455 -338 1521 -322
rect 1569 -326 1599 -300
rect 1665 -322 1695 -300
rect 1455 -372 1471 -338
rect 1505 -372 1521 -338
rect 1455 -388 1521 -372
rect 1647 -338 1713 -322
rect 1761 -326 1791 -300
rect 1857 -322 1887 -300
rect 1647 -372 1663 -338
rect 1697 -372 1713 -338
rect 1647 -388 1713 -372
rect 1839 -338 1905 -322
rect 1953 -326 1983 -300
rect 1839 -372 1855 -338
rect 1889 -372 1905 -338
rect 1839 -388 1905 -372
<< polycont >>
rect -1889 338 -1855 372
rect -1697 338 -1663 372
rect -1505 338 -1471 372
rect -1313 338 -1279 372
rect -1121 338 -1087 372
rect -929 338 -895 372
rect -737 338 -703 372
rect -545 338 -511 372
rect -353 338 -319 372
rect -161 338 -127 372
rect 31 338 65 372
rect 223 338 257 372
rect 415 338 449 372
rect 607 338 641 372
rect 799 338 833 372
rect 991 338 1025 372
rect 1183 338 1217 372
rect 1375 338 1409 372
rect 1567 338 1601 372
rect 1759 338 1793 372
rect 1951 338 1985 372
rect -1985 -372 -1951 -338
rect -1793 -372 -1759 -338
rect -1601 -372 -1567 -338
rect -1409 -372 -1375 -338
rect -1217 -372 -1183 -338
rect -1025 -372 -991 -338
rect -833 -372 -799 -338
rect -641 -372 -607 -338
rect -449 -372 -415 -338
rect -257 -372 -223 -338
rect -65 -372 -31 -338
rect 127 -372 161 -338
rect 319 -372 353 -338
rect 511 -372 545 -338
rect 703 -372 737 -338
rect 895 -372 929 -338
rect 1087 -372 1121 -338
rect 1279 -372 1313 -338
rect 1471 -372 1505 -338
rect 1663 -372 1697 -338
rect 1855 -372 1889 -338
<< locali >>
rect -2147 440 -2051 474
rect 2051 440 2147 474
rect -2147 378 -2113 440
rect 2113 378 2147 440
rect -1905 338 -1889 372
rect -1855 338 -1839 372
rect -1713 338 -1697 372
rect -1663 338 -1647 372
rect -1521 338 -1505 372
rect -1471 338 -1455 372
rect -1329 338 -1313 372
rect -1279 338 -1263 372
rect -1137 338 -1121 372
rect -1087 338 -1071 372
rect -945 338 -929 372
rect -895 338 -879 372
rect -753 338 -737 372
rect -703 338 -687 372
rect -561 338 -545 372
rect -511 338 -495 372
rect -369 338 -353 372
rect -319 338 -303 372
rect -177 338 -161 372
rect -127 338 -111 372
rect 15 338 31 372
rect 65 338 81 372
rect 207 338 223 372
rect 257 338 273 372
rect 399 338 415 372
rect 449 338 465 372
rect 591 338 607 372
rect 641 338 657 372
rect 783 338 799 372
rect 833 338 849 372
rect 975 338 991 372
rect 1025 338 1041 372
rect 1167 338 1183 372
rect 1217 338 1233 372
rect 1359 338 1375 372
rect 1409 338 1425 372
rect 1551 338 1567 372
rect 1601 338 1617 372
rect 1743 338 1759 372
rect 1793 338 1809 372
rect 1935 338 1951 372
rect 1985 338 2001 372
rect -2033 288 -1999 304
rect -2033 -304 -1999 -288
rect -1937 288 -1903 304
rect -1937 -304 -1903 -288
rect -1841 288 -1807 304
rect -1841 -304 -1807 -288
rect -1745 288 -1711 304
rect -1745 -304 -1711 -288
rect -1649 288 -1615 304
rect -1649 -304 -1615 -288
rect -1553 288 -1519 304
rect -1553 -304 -1519 -288
rect -1457 288 -1423 304
rect -1457 -304 -1423 -288
rect -1361 288 -1327 304
rect -1361 -304 -1327 -288
rect -1265 288 -1231 304
rect -1265 -304 -1231 -288
rect -1169 288 -1135 304
rect -1169 -304 -1135 -288
rect -1073 288 -1039 304
rect -1073 -304 -1039 -288
rect -977 288 -943 304
rect -977 -304 -943 -288
rect -881 288 -847 304
rect -881 -304 -847 -288
rect -785 288 -751 304
rect -785 -304 -751 -288
rect -689 288 -655 304
rect -689 -304 -655 -288
rect -593 288 -559 304
rect -593 -304 -559 -288
rect -497 288 -463 304
rect -497 -304 -463 -288
rect -401 288 -367 304
rect -401 -304 -367 -288
rect -305 288 -271 304
rect -305 -304 -271 -288
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect 271 288 305 304
rect 271 -304 305 -288
rect 367 288 401 304
rect 367 -304 401 -288
rect 463 288 497 304
rect 463 -304 497 -288
rect 559 288 593 304
rect 559 -304 593 -288
rect 655 288 689 304
rect 655 -304 689 -288
rect 751 288 785 304
rect 751 -304 785 -288
rect 847 288 881 304
rect 847 -304 881 -288
rect 943 288 977 304
rect 943 -304 977 -288
rect 1039 288 1073 304
rect 1039 -304 1073 -288
rect 1135 288 1169 304
rect 1135 -304 1169 -288
rect 1231 288 1265 304
rect 1231 -304 1265 -288
rect 1327 288 1361 304
rect 1327 -304 1361 -288
rect 1423 288 1457 304
rect 1423 -304 1457 -288
rect 1519 288 1553 304
rect 1519 -304 1553 -288
rect 1615 288 1649 304
rect 1615 -304 1649 -288
rect 1711 288 1745 304
rect 1711 -304 1745 -288
rect 1807 288 1841 304
rect 1807 -304 1841 -288
rect 1903 288 1937 304
rect 1903 -304 1937 -288
rect 1999 288 2033 304
rect 1999 -304 2033 -288
rect -2001 -372 -1985 -338
rect -1951 -372 -1935 -338
rect -1809 -372 -1793 -338
rect -1759 -372 -1743 -338
rect -1617 -372 -1601 -338
rect -1567 -372 -1551 -338
rect -1425 -372 -1409 -338
rect -1375 -372 -1359 -338
rect -1233 -372 -1217 -338
rect -1183 -372 -1167 -338
rect -1041 -372 -1025 -338
rect -991 -372 -975 -338
rect -849 -372 -833 -338
rect -799 -372 -783 -338
rect -657 -372 -641 -338
rect -607 -372 -591 -338
rect -465 -372 -449 -338
rect -415 -372 -399 -338
rect -273 -372 -257 -338
rect -223 -372 -207 -338
rect -81 -372 -65 -338
rect -31 -372 -15 -338
rect 111 -372 127 -338
rect 161 -372 177 -338
rect 303 -372 319 -338
rect 353 -372 369 -338
rect 495 -372 511 -338
rect 545 -372 561 -338
rect 687 -372 703 -338
rect 737 -372 753 -338
rect 879 -372 895 -338
rect 929 -372 945 -338
rect 1071 -372 1087 -338
rect 1121 -372 1137 -338
rect 1263 -372 1279 -338
rect 1313 -372 1329 -338
rect 1455 -372 1471 -338
rect 1505 -372 1521 -338
rect 1647 -372 1663 -338
rect 1697 -372 1713 -338
rect 1839 -372 1855 -338
rect 1889 -372 1905 -338
rect -2147 -440 -2113 -378
rect 2113 -440 2147 -378
rect -2147 -474 -2051 -440
rect 2051 -474 2147 -440
<< viali >>
rect -1889 338 -1855 372
rect -1697 338 -1663 372
rect -1505 338 -1471 372
rect -1313 338 -1279 372
rect -1121 338 -1087 372
rect -929 338 -895 372
rect -737 338 -703 372
rect -545 338 -511 372
rect -353 338 -319 372
rect -161 338 -127 372
rect 31 338 65 372
rect 223 338 257 372
rect 415 338 449 372
rect 607 338 641 372
rect 799 338 833 372
rect 991 338 1025 372
rect 1183 338 1217 372
rect 1375 338 1409 372
rect 1567 338 1601 372
rect 1759 338 1793 372
rect 1951 338 1985 372
rect -2033 -288 -1999 288
rect -1937 -288 -1903 288
rect -1841 -288 -1807 288
rect -1745 -288 -1711 288
rect -1649 -288 -1615 288
rect -1553 -288 -1519 288
rect -1457 -288 -1423 288
rect -1361 -288 -1327 288
rect -1265 -288 -1231 288
rect -1169 -288 -1135 288
rect -1073 -288 -1039 288
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
rect 1039 -288 1073 288
rect 1135 -288 1169 288
rect 1231 -288 1265 288
rect 1327 -288 1361 288
rect 1423 -288 1457 288
rect 1519 -288 1553 288
rect 1615 -288 1649 288
rect 1711 -288 1745 288
rect 1807 -288 1841 288
rect 1903 -288 1937 288
rect 1999 -288 2033 288
rect -1985 -372 -1951 -338
rect -1793 -372 -1759 -338
rect -1601 -372 -1567 -338
rect -1409 -372 -1375 -338
rect -1217 -372 -1183 -338
rect -1025 -372 -991 -338
rect -833 -372 -799 -338
rect -641 -372 -607 -338
rect -449 -372 -415 -338
rect -257 -372 -223 -338
rect -65 -372 -31 -338
rect 127 -372 161 -338
rect 319 -372 353 -338
rect 511 -372 545 -338
rect 703 -372 737 -338
rect 895 -372 929 -338
rect 1087 -372 1121 -338
rect 1279 -372 1313 -338
rect 1471 -372 1505 -338
rect 1663 -372 1697 -338
rect 1855 -372 1889 -338
<< metal1 >>
rect -1901 372 -1843 378
rect -1901 338 -1889 372
rect -1855 338 -1843 372
rect -1901 332 -1843 338
rect -1709 372 -1651 378
rect -1709 338 -1697 372
rect -1663 338 -1651 372
rect -1709 332 -1651 338
rect -1517 372 -1459 378
rect -1517 338 -1505 372
rect -1471 338 -1459 372
rect -1517 332 -1459 338
rect -1325 372 -1267 378
rect -1325 338 -1313 372
rect -1279 338 -1267 372
rect -1325 332 -1267 338
rect -1133 372 -1075 378
rect -1133 338 -1121 372
rect -1087 338 -1075 372
rect -1133 332 -1075 338
rect -941 372 -883 378
rect -941 338 -929 372
rect -895 338 -883 372
rect -941 332 -883 338
rect -749 372 -691 378
rect -749 338 -737 372
rect -703 338 -691 372
rect -749 332 -691 338
rect -557 372 -499 378
rect -557 338 -545 372
rect -511 338 -499 372
rect -557 332 -499 338
rect -365 372 -307 378
rect -365 338 -353 372
rect -319 338 -307 372
rect -365 332 -307 338
rect -173 372 -115 378
rect -173 338 -161 372
rect -127 338 -115 372
rect -173 332 -115 338
rect 19 372 77 378
rect 19 338 31 372
rect 65 338 77 372
rect 19 332 77 338
rect 211 372 269 378
rect 211 338 223 372
rect 257 338 269 372
rect 211 332 269 338
rect 403 372 461 378
rect 403 338 415 372
rect 449 338 461 372
rect 403 332 461 338
rect 595 372 653 378
rect 595 338 607 372
rect 641 338 653 372
rect 595 332 653 338
rect 787 372 845 378
rect 787 338 799 372
rect 833 338 845 372
rect 787 332 845 338
rect 979 372 1037 378
rect 979 338 991 372
rect 1025 338 1037 372
rect 979 332 1037 338
rect 1171 372 1229 378
rect 1171 338 1183 372
rect 1217 338 1229 372
rect 1171 332 1229 338
rect 1363 372 1421 378
rect 1363 338 1375 372
rect 1409 338 1421 372
rect 1363 332 1421 338
rect 1555 372 1613 378
rect 1555 338 1567 372
rect 1601 338 1613 372
rect 1555 332 1613 338
rect 1747 372 1805 378
rect 1747 338 1759 372
rect 1793 338 1805 372
rect 1747 332 1805 338
rect 1939 372 1997 378
rect 1939 338 1951 372
rect 1985 338 1997 372
rect 1939 332 1997 338
rect -2039 288 -1993 300
rect -2039 -288 -2033 288
rect -1999 -288 -1993 288
rect -2039 -300 -1993 -288
rect -1943 288 -1897 300
rect -1943 -288 -1937 288
rect -1903 -288 -1897 288
rect -1943 -300 -1897 -288
rect -1847 288 -1801 300
rect -1847 -288 -1841 288
rect -1807 -288 -1801 288
rect -1847 -300 -1801 -288
rect -1751 288 -1705 300
rect -1751 -288 -1745 288
rect -1711 -288 -1705 288
rect -1751 -300 -1705 -288
rect -1655 288 -1609 300
rect -1655 -288 -1649 288
rect -1615 -288 -1609 288
rect -1655 -300 -1609 -288
rect -1559 288 -1513 300
rect -1559 -288 -1553 288
rect -1519 -288 -1513 288
rect -1559 -300 -1513 -288
rect -1463 288 -1417 300
rect -1463 -288 -1457 288
rect -1423 -288 -1417 288
rect -1463 -300 -1417 -288
rect -1367 288 -1321 300
rect -1367 -288 -1361 288
rect -1327 -288 -1321 288
rect -1367 -300 -1321 -288
rect -1271 288 -1225 300
rect -1271 -288 -1265 288
rect -1231 -288 -1225 288
rect -1271 -300 -1225 -288
rect -1175 288 -1129 300
rect -1175 -288 -1169 288
rect -1135 -288 -1129 288
rect -1175 -300 -1129 -288
rect -1079 288 -1033 300
rect -1079 -288 -1073 288
rect -1039 -288 -1033 288
rect -1079 -300 -1033 -288
rect -983 288 -937 300
rect -983 -288 -977 288
rect -943 -288 -937 288
rect -983 -300 -937 -288
rect -887 288 -841 300
rect -887 -288 -881 288
rect -847 -288 -841 288
rect -887 -300 -841 -288
rect -791 288 -745 300
rect -791 -288 -785 288
rect -751 -288 -745 288
rect -791 -300 -745 -288
rect -695 288 -649 300
rect -695 -288 -689 288
rect -655 -288 -649 288
rect -695 -300 -649 -288
rect -599 288 -553 300
rect -599 -288 -593 288
rect -559 -288 -553 288
rect -599 -300 -553 -288
rect -503 288 -457 300
rect -503 -288 -497 288
rect -463 -288 -457 288
rect -503 -300 -457 -288
rect -407 288 -361 300
rect -407 -288 -401 288
rect -367 -288 -361 288
rect -407 -300 -361 -288
rect -311 288 -265 300
rect -311 -288 -305 288
rect -271 -288 -265 288
rect -311 -300 -265 -288
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect 265 288 311 300
rect 265 -288 271 288
rect 305 -288 311 288
rect 265 -300 311 -288
rect 361 288 407 300
rect 361 -288 367 288
rect 401 -288 407 288
rect 361 -300 407 -288
rect 457 288 503 300
rect 457 -288 463 288
rect 497 -288 503 288
rect 457 -300 503 -288
rect 553 288 599 300
rect 553 -288 559 288
rect 593 -288 599 288
rect 553 -300 599 -288
rect 649 288 695 300
rect 649 -288 655 288
rect 689 -288 695 288
rect 649 -300 695 -288
rect 745 288 791 300
rect 745 -288 751 288
rect 785 -288 791 288
rect 745 -300 791 -288
rect 841 288 887 300
rect 841 -288 847 288
rect 881 -288 887 288
rect 841 -300 887 -288
rect 937 288 983 300
rect 937 -288 943 288
rect 977 -288 983 288
rect 937 -300 983 -288
rect 1033 288 1079 300
rect 1033 -288 1039 288
rect 1073 -288 1079 288
rect 1033 -300 1079 -288
rect 1129 288 1175 300
rect 1129 -288 1135 288
rect 1169 -288 1175 288
rect 1129 -300 1175 -288
rect 1225 288 1271 300
rect 1225 -288 1231 288
rect 1265 -288 1271 288
rect 1225 -300 1271 -288
rect 1321 288 1367 300
rect 1321 -288 1327 288
rect 1361 -288 1367 288
rect 1321 -300 1367 -288
rect 1417 288 1463 300
rect 1417 -288 1423 288
rect 1457 -288 1463 288
rect 1417 -300 1463 -288
rect 1513 288 1559 300
rect 1513 -288 1519 288
rect 1553 -288 1559 288
rect 1513 -300 1559 -288
rect 1609 288 1655 300
rect 1609 -288 1615 288
rect 1649 -288 1655 288
rect 1609 -300 1655 -288
rect 1705 288 1751 300
rect 1705 -288 1711 288
rect 1745 -288 1751 288
rect 1705 -300 1751 -288
rect 1801 288 1847 300
rect 1801 -288 1807 288
rect 1841 -288 1847 288
rect 1801 -300 1847 -288
rect 1897 288 1943 300
rect 1897 -288 1903 288
rect 1937 -288 1943 288
rect 1897 -300 1943 -288
rect 1993 288 2039 300
rect 1993 -288 1999 288
rect 2033 -288 2039 288
rect 1993 -300 2039 -288
rect -1997 -338 -1939 -332
rect -1997 -372 -1985 -338
rect -1951 -372 -1939 -338
rect -1997 -378 -1939 -372
rect -1805 -338 -1747 -332
rect -1805 -372 -1793 -338
rect -1759 -372 -1747 -338
rect -1805 -378 -1747 -372
rect -1613 -338 -1555 -332
rect -1613 -372 -1601 -338
rect -1567 -372 -1555 -338
rect -1613 -378 -1555 -372
rect -1421 -338 -1363 -332
rect -1421 -372 -1409 -338
rect -1375 -372 -1363 -338
rect -1421 -378 -1363 -372
rect -1229 -338 -1171 -332
rect -1229 -372 -1217 -338
rect -1183 -372 -1171 -338
rect -1229 -378 -1171 -372
rect -1037 -338 -979 -332
rect -1037 -372 -1025 -338
rect -991 -372 -979 -338
rect -1037 -378 -979 -372
rect -845 -338 -787 -332
rect -845 -372 -833 -338
rect -799 -372 -787 -338
rect -845 -378 -787 -372
rect -653 -338 -595 -332
rect -653 -372 -641 -338
rect -607 -372 -595 -338
rect -653 -378 -595 -372
rect -461 -338 -403 -332
rect -461 -372 -449 -338
rect -415 -372 -403 -338
rect -461 -378 -403 -372
rect -269 -338 -211 -332
rect -269 -372 -257 -338
rect -223 -372 -211 -338
rect -269 -378 -211 -372
rect -77 -338 -19 -332
rect -77 -372 -65 -338
rect -31 -372 -19 -338
rect -77 -378 -19 -372
rect 115 -338 173 -332
rect 115 -372 127 -338
rect 161 -372 173 -338
rect 115 -378 173 -372
rect 307 -338 365 -332
rect 307 -372 319 -338
rect 353 -372 365 -338
rect 307 -378 365 -372
rect 499 -338 557 -332
rect 499 -372 511 -338
rect 545 -372 557 -338
rect 499 -378 557 -372
rect 691 -338 749 -332
rect 691 -372 703 -338
rect 737 -372 749 -338
rect 691 -378 749 -372
rect 883 -338 941 -332
rect 883 -372 895 -338
rect 929 -372 941 -338
rect 883 -378 941 -372
rect 1075 -338 1133 -332
rect 1075 -372 1087 -338
rect 1121 -372 1133 -338
rect 1075 -378 1133 -372
rect 1267 -338 1325 -332
rect 1267 -372 1279 -338
rect 1313 -372 1325 -338
rect 1267 -378 1325 -372
rect 1459 -338 1517 -332
rect 1459 -372 1471 -338
rect 1505 -372 1517 -338
rect 1459 -378 1517 -372
rect 1651 -338 1709 -332
rect 1651 -372 1663 -338
rect 1697 -372 1709 -338
rect 1651 -378 1709 -372
rect 1843 -338 1901 -332
rect 1843 -372 1855 -338
rect 1889 -372 1901 -338
rect 1843 -378 1901 -372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -2130 -457 2130 457
string parameters w 3 l 0.150 m 1 nf 42 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
