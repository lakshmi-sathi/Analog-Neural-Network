magic
tech sky130A
magscale 1 2
timestamp 1627805856
<< xpolycontact >>
rect -35 77 35 509
rect -35 -509 35 -77
<< xpolyres >>
rect -35 -77 35 77
<< viali >>
rect -19 94 19 491
rect -19 -491 19 -94
<< metal1 >>
rect -25 491 25 503
rect -25 94 -19 491
rect 19 94 25 491
rect -25 82 25 94
rect -25 -94 25 -82
rect -25 -491 -19 -94
rect 19 -491 25 -94
rect -25 -503 25 -491
<< res0p35 >>
rect -37 -79 37 79
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 0.77 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.085k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
