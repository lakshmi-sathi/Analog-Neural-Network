magic
tech sky130A
magscale 1 2
timestamp 1628080314
<< error_p >>
rect -269 511 -211 517
rect -77 511 -19 517
rect 115 511 173 517
rect 307 511 365 517
rect -269 477 -257 511
rect -77 477 -65 511
rect 115 477 127 511
rect 307 477 319 511
rect -269 471 -211 477
rect -77 471 -19 477
rect 115 471 173 477
rect 307 471 365 477
rect -365 -477 -307 -471
rect -173 -477 -115 -471
rect 19 -477 77 -471
rect 211 -477 269 -471
rect -365 -511 -353 -477
rect -173 -511 -161 -477
rect 19 -511 31 -477
rect 211 -511 223 -477
rect -365 -517 -307 -511
rect -173 -517 -115 -511
rect 19 -517 77 -511
rect 211 -517 269 -511
<< nwell >>
rect -551 -649 551 649
<< pmos >>
rect -351 -430 -321 430
rect -255 -430 -225 430
rect -159 -430 -129 430
rect -63 -430 -33 430
rect 33 -430 63 430
rect 129 -430 159 430
rect 225 -430 255 430
rect 321 -430 351 430
<< pdiff >>
rect -413 418 -351 430
rect -413 -418 -401 418
rect -367 -418 -351 418
rect -413 -430 -351 -418
rect -321 418 -255 430
rect -321 -418 -305 418
rect -271 -418 -255 418
rect -321 -430 -255 -418
rect -225 418 -159 430
rect -225 -418 -209 418
rect -175 -418 -159 418
rect -225 -430 -159 -418
rect -129 418 -63 430
rect -129 -418 -113 418
rect -79 -418 -63 418
rect -129 -430 -63 -418
rect -33 418 33 430
rect -33 -418 -17 418
rect 17 -418 33 418
rect -33 -430 33 -418
rect 63 418 129 430
rect 63 -418 79 418
rect 113 -418 129 418
rect 63 -430 129 -418
rect 159 418 225 430
rect 159 -418 175 418
rect 209 -418 225 418
rect 159 -430 225 -418
rect 255 418 321 430
rect 255 -418 271 418
rect 305 -418 321 418
rect 255 -430 321 -418
rect 351 418 413 430
rect 351 -418 367 418
rect 401 -418 413 418
rect 351 -430 413 -418
<< pdiffc >>
rect -401 -418 -367 418
rect -305 -418 -271 418
rect -209 -418 -175 418
rect -113 -418 -79 418
rect -17 -418 17 418
rect 79 -418 113 418
rect 175 -418 209 418
rect 271 -418 305 418
rect 367 -418 401 418
<< nsubdiff >>
rect -515 579 -419 613
rect 419 579 515 613
rect -515 517 -481 579
rect 481 517 515 579
rect -515 -579 -481 -517
rect 481 -579 515 -517
rect -515 -613 -419 -579
rect 419 -613 515 -579
<< nsubdiffcont >>
rect -419 579 419 613
rect -515 -517 -481 517
rect 481 -517 515 517
rect -419 -613 419 -579
<< poly >>
rect -273 511 -207 527
rect -273 477 -257 511
rect -223 477 -207 511
rect -273 461 -207 477
rect -81 511 -15 527
rect -81 477 -65 511
rect -31 477 -15 511
rect -81 461 -15 477
rect 111 511 177 527
rect 111 477 127 511
rect 161 477 177 511
rect 111 461 177 477
rect 303 511 369 527
rect 303 477 319 511
rect 353 477 369 511
rect 303 461 369 477
rect -351 430 -321 456
rect -255 430 -225 461
rect -159 430 -129 456
rect -63 430 -33 461
rect 33 430 63 456
rect 129 430 159 461
rect 225 430 255 456
rect 321 430 351 461
rect -351 -461 -321 -430
rect -255 -456 -225 -430
rect -159 -461 -129 -430
rect -63 -456 -33 -430
rect 33 -461 63 -430
rect 129 -456 159 -430
rect 225 -461 255 -430
rect 321 -456 351 -430
rect -369 -477 -303 -461
rect -369 -511 -353 -477
rect -319 -511 -303 -477
rect -369 -527 -303 -511
rect -177 -477 -111 -461
rect -177 -511 -161 -477
rect -127 -511 -111 -477
rect -177 -527 -111 -511
rect 15 -477 81 -461
rect 15 -511 31 -477
rect 65 -511 81 -477
rect 15 -527 81 -511
rect 207 -477 273 -461
rect 207 -511 223 -477
rect 257 -511 273 -477
rect 207 -527 273 -511
<< polycont >>
rect -257 477 -223 511
rect -65 477 -31 511
rect 127 477 161 511
rect 319 477 353 511
rect -353 -511 -319 -477
rect -161 -511 -127 -477
rect 31 -511 65 -477
rect 223 -511 257 -477
<< locali >>
rect -515 579 -419 613
rect 419 579 515 613
rect -515 517 -481 579
rect 481 517 515 579
rect -273 477 -257 511
rect -223 477 -207 511
rect -81 477 -65 511
rect -31 477 -15 511
rect 111 477 127 511
rect 161 477 177 511
rect 303 477 319 511
rect 353 477 369 511
rect -401 418 -367 434
rect -401 -434 -367 -418
rect -305 418 -271 434
rect -305 -434 -271 -418
rect -209 418 -175 434
rect -209 -434 -175 -418
rect -113 418 -79 434
rect -113 -434 -79 -418
rect -17 418 17 434
rect -17 -434 17 -418
rect 79 418 113 434
rect 79 -434 113 -418
rect 175 418 209 434
rect 175 -434 209 -418
rect 271 418 305 434
rect 271 -434 305 -418
rect 367 418 401 434
rect 367 -434 401 -418
rect -369 -511 -353 -477
rect -319 -511 -303 -477
rect -177 -511 -161 -477
rect -127 -511 -111 -477
rect 15 -511 31 -477
rect 65 -511 81 -477
rect 207 -511 223 -477
rect 257 -511 273 -477
rect -515 -579 -481 -517
rect 481 -579 515 -517
rect -515 -613 -419 -579
rect 419 -613 515 -579
<< viali >>
rect -257 477 -223 511
rect -65 477 -31 511
rect 127 477 161 511
rect 319 477 353 511
rect -401 -418 -367 418
rect -305 -418 -271 418
rect -209 -418 -175 418
rect -113 -418 -79 418
rect -17 -418 17 418
rect 79 -418 113 418
rect 175 -418 209 418
rect 271 -418 305 418
rect 367 -418 401 418
rect -353 -511 -319 -477
rect -161 -511 -127 -477
rect 31 -511 65 -477
rect 223 -511 257 -477
<< metal1 >>
rect -269 511 -211 517
rect -269 477 -257 511
rect -223 477 -211 511
rect -269 471 -211 477
rect -77 511 -19 517
rect -77 477 -65 511
rect -31 477 -19 511
rect -77 471 -19 477
rect 115 511 173 517
rect 115 477 127 511
rect 161 477 173 511
rect 115 471 173 477
rect 307 511 365 517
rect 307 477 319 511
rect 353 477 365 511
rect 307 471 365 477
rect -407 418 -361 430
rect -407 -418 -401 418
rect -367 -418 -361 418
rect -407 -430 -361 -418
rect -311 418 -265 430
rect -311 -418 -305 418
rect -271 -418 -265 418
rect -311 -430 -265 -418
rect -215 418 -169 430
rect -215 -418 -209 418
rect -175 -418 -169 418
rect -215 -430 -169 -418
rect -119 418 -73 430
rect -119 -418 -113 418
rect -79 -418 -73 418
rect -119 -430 -73 -418
rect -23 418 23 430
rect -23 -418 -17 418
rect 17 -418 23 418
rect -23 -430 23 -418
rect 73 418 119 430
rect 73 -418 79 418
rect 113 -418 119 418
rect 73 -430 119 -418
rect 169 418 215 430
rect 169 -418 175 418
rect 209 -418 215 418
rect 169 -430 215 -418
rect 265 418 311 430
rect 265 -418 271 418
rect 305 -418 311 418
rect 265 -430 311 -418
rect 361 418 407 430
rect 361 -418 367 418
rect 401 -418 407 418
rect 361 -430 407 -418
rect -365 -477 -307 -471
rect -365 -511 -353 -477
rect -319 -511 -307 -477
rect -365 -517 -307 -511
rect -173 -477 -115 -471
rect -173 -511 -161 -477
rect -127 -511 -115 -477
rect -173 -517 -115 -511
rect 19 -477 77 -471
rect 19 -511 31 -477
rect 65 -511 77 -477
rect 19 -517 77 -511
rect 211 -477 269 -471
rect 211 -511 223 -477
rect 257 -511 269 -477
rect 211 -517 269 -511
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -498 -596 498 596
string parameters w 4.3 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
