magic
tech sky130A
magscale 1 2
timestamp 1627922418
<< pwell >>
rect -201 -981 201 981
<< psubdiff >>
rect -165 911 -69 945
rect 69 911 165 945
rect -165 849 -131 911
rect 131 849 165 911
rect -165 -911 -131 -849
rect 131 -911 165 -849
rect -165 -945 -69 -911
rect 69 -945 165 -911
<< psubdiffcont >>
rect -69 911 69 945
rect -165 -849 -131 849
rect 131 -849 165 849
rect -69 -945 69 -911
<< xpolycontact >>
rect -35 383 35 815
rect -35 -815 35 -383
<< xpolyres >>
rect -35 -383 35 383
<< locali >>
rect -165 911 -69 945
rect 69 911 165 945
rect -165 849 -131 911
rect 131 849 165 911
rect -165 -911 -131 -849
rect 131 -911 165 -849
rect -165 -945 -69 -911
rect 69 -945 165 -911
<< viali >>
rect -19 400 19 797
rect -19 -797 19 -400
<< metal1 >>
rect -25 797 25 809
rect -25 400 -19 797
rect 19 400 25 797
rect -25 388 25 400
rect -25 -400 25 -388
rect -25 -797 -19 -400
rect 19 -797 25 -400
rect -25 -809 25 -797
<< res0p35 >>
rect -37 -385 37 385
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string FIXED_BBOX -148 -928 148 928
string parameters w 0.350 l 3.83 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 22.571k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
