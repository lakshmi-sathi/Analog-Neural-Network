magic
tech sky130A
magscale 1 2
timestamp 1628080314
<< error_p >>
rect 19 582 77 588
rect 19 548 31 582
rect 19 542 77 548
rect -77 -548 -19 -542
rect -77 -582 -65 -548
rect -77 -588 -19 -582
<< pwell >>
rect -263 -720 263 720
<< nmos >>
rect -63 -510 -33 510
rect 33 -510 63 510
<< ndiff >>
rect -125 498 -63 510
rect -125 -498 -113 498
rect -79 -498 -63 498
rect -125 -510 -63 -498
rect -33 498 33 510
rect -33 -498 -17 498
rect 17 -498 33 498
rect -33 -510 33 -498
rect 63 498 125 510
rect 63 -498 79 498
rect 113 -498 125 498
rect 63 -510 125 -498
<< ndiffc >>
rect -113 -498 -79 498
rect -17 -498 17 498
rect 79 -498 113 498
<< psubdiff >>
rect -227 650 -131 684
rect 131 650 227 684
rect -227 588 -193 650
rect 193 588 227 650
rect -227 -650 -193 -588
rect 193 -650 227 -588
rect -227 -684 -131 -650
rect 131 -684 227 -650
<< psubdiffcont >>
rect -131 650 131 684
rect -227 -588 -193 588
rect 193 -588 227 588
rect -131 -684 131 -650
<< poly >>
rect 15 582 81 598
rect 15 548 31 582
rect 65 548 81 582
rect -63 510 -33 536
rect 15 532 81 548
rect 33 510 63 532
rect -63 -532 -33 -510
rect -81 -548 -15 -532
rect 33 -536 63 -510
rect -81 -582 -65 -548
rect -31 -582 -15 -548
rect -81 -598 -15 -582
<< polycont >>
rect 31 548 65 582
rect -65 -582 -31 -548
<< locali >>
rect -227 650 -131 684
rect 131 650 227 684
rect -227 588 -193 650
rect 193 588 227 650
rect 15 548 31 582
rect 65 548 81 582
rect -113 498 -79 514
rect -113 -514 -79 -498
rect -17 498 17 514
rect -17 -514 17 -498
rect 79 498 113 514
rect 79 -514 113 -498
rect -81 -582 -65 -548
rect -31 -582 -15 -548
rect -227 -650 -193 -588
rect 193 -650 227 -588
rect -227 -684 -131 -650
rect 131 -684 227 -650
<< viali >>
rect 31 548 65 582
rect -113 -498 -79 498
rect -17 -498 17 498
rect 79 -498 113 498
rect -65 -582 -31 -548
<< metal1 >>
rect 19 582 77 588
rect 19 548 31 582
rect 65 548 77 582
rect 19 542 77 548
rect -119 498 -73 510
rect -119 -498 -113 498
rect -79 -498 -73 498
rect -119 -510 -73 -498
rect -23 498 23 510
rect -23 -498 -17 498
rect 17 -498 23 498
rect -23 -510 23 -498
rect 73 498 119 510
rect 73 -498 79 498
rect 113 -498 119 498
rect 73 -510 119 -498
rect -77 -548 -19 -542
rect -77 -582 -65 -548
rect -31 -582 -19 -548
rect -77 -588 -19 -582
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -210 -667 210 667
string parameters w 5.1 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
