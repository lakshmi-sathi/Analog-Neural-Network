magic
tech sky130A
magscale 1 2
timestamp 1627032624
<< xpolycontact >>
rect -35 536 35 968
rect -35 -968 35 -536
<< ppolyres >>
rect -35 -536 35 536
<< viali >>
rect -19 553 19 950
rect -19 -950 19 -553
<< metal1 >>
rect -25 950 25 962
rect -25 553 -19 950
rect 19 553 25 950
rect -25 541 25 553
rect -25 -553 25 -541
rect -25 -950 -19 -553
rect 19 -950 25 -553
rect -25 -962 25 -950
<< res0p35 >>
rect -37 -538 37 538
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string parameters w 0.350 l 5.36 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 5.007k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 0.350 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
