magic
tech sky130A
magscale 1 2
timestamp 1628058135
<< error_p >>
rect -29 1001 29 1007
rect -29 967 -17 1001
rect -29 961 29 967
<< pwell >>
rect -211 -1139 211 1139
<< nmos >>
rect -15 -991 15 929
<< ndiff >>
rect -73 917 -15 929
rect -73 -979 -61 917
rect -27 -979 -15 917
rect -73 -991 -15 -979
rect 15 917 73 929
rect 15 -979 27 917
rect 61 -979 73 917
rect 15 -991 73 -979
<< ndiffc >>
rect -61 -979 -27 917
rect 27 -979 61 917
<< psubdiff >>
rect -175 1069 -79 1103
rect 79 1069 175 1103
rect -175 1007 -141 1069
rect 141 1007 175 1069
rect -175 -1069 -141 -1007
rect 141 -1069 175 -1007
rect -175 -1103 -79 -1069
rect 79 -1103 175 -1069
<< psubdiffcont >>
rect -79 1069 79 1103
rect -175 -1007 -141 1007
rect 141 -1007 175 1007
rect -79 -1103 79 -1069
<< poly >>
rect -33 1001 33 1017
rect -33 967 -17 1001
rect 17 967 33 1001
rect -33 951 33 967
rect -15 929 15 951
rect -15 -1017 15 -991
<< polycont >>
rect -17 967 17 1001
<< locali >>
rect -175 1069 -79 1103
rect 79 1069 175 1103
rect -175 1007 -141 1069
rect 141 1007 175 1069
rect -33 967 -17 1001
rect 17 967 33 1001
rect -61 917 -27 933
rect -61 -995 -27 -979
rect 27 917 61 933
rect 27 -995 61 -979
rect -175 -1069 -141 -1007
rect 141 -1069 175 -1007
rect -175 -1103 -79 -1069
rect 79 -1103 175 -1069
<< viali >>
rect -17 967 17 1001
rect -61 -979 -27 917
rect 27 -979 61 917
<< metal1 >>
rect -29 1001 29 1007
rect -29 967 -17 1001
rect 17 967 29 1001
rect -29 961 29 967
rect -67 917 -21 929
rect -67 -979 -61 917
rect -27 -979 -21 917
rect -67 -991 -21 -979
rect 21 917 67 929
rect 21 -979 27 917
rect 61 -979 67 917
rect 21 -991 67 -979
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -1086 158 1086
string parameters w 9.6 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
