magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_p >>
rect -845 373 -787 379
rect -653 373 -595 379
rect -461 373 -403 379
rect -269 373 -211 379
rect -77 373 -19 379
rect 115 373 173 379
rect 307 373 365 379
rect 499 373 557 379
rect 691 373 749 379
rect -845 339 -833 373
rect -653 339 -641 373
rect -461 339 -449 373
rect -269 339 -257 373
rect -77 339 -65 373
rect 115 339 127 373
rect 307 339 319 373
rect 499 339 511 373
rect 691 339 703 373
rect -845 333 -787 339
rect -653 333 -595 339
rect -461 333 -403 339
rect -269 333 -211 339
rect -77 333 -19 339
rect 115 333 173 339
rect 307 333 365 339
rect 499 333 557 339
rect 691 333 749 339
rect -749 71 -691 77
rect -557 71 -499 77
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect 595 71 653 77
rect 787 71 845 77
rect -749 37 -737 71
rect -557 37 -545 71
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect 595 37 607 71
rect 787 37 799 71
rect -749 31 -691 37
rect -557 31 -499 37
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect 595 31 653 37
rect 787 31 845 37
rect -749 -37 -691 -31
rect -557 -37 -499 -31
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect 595 -37 653 -31
rect 787 -37 845 -31
rect -749 -71 -737 -37
rect -557 -71 -545 -37
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect 595 -71 607 -37
rect 787 -71 799 -37
rect -749 -77 -691 -71
rect -557 -77 -499 -71
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect 595 -77 653 -71
rect 787 -77 845 -71
rect -845 -339 -787 -333
rect -653 -339 -595 -333
rect -461 -339 -403 -333
rect -269 -339 -211 -333
rect -77 -339 -19 -333
rect 115 -339 173 -333
rect 307 -339 365 -333
rect 499 -339 557 -333
rect 691 -339 749 -333
rect -845 -373 -833 -339
rect -653 -373 -641 -339
rect -461 -373 -449 -339
rect -269 -373 -257 -339
rect -77 -373 -65 -339
rect 115 -373 127 -339
rect 307 -373 319 -339
rect 499 -373 511 -339
rect 691 -373 703 -339
rect -845 -379 -787 -373
rect -653 -379 -595 -373
rect -461 -379 -403 -373
rect -269 -379 -211 -373
rect -77 -379 -19 -373
rect 115 -379 173 -373
rect 307 -379 365 -373
rect 499 -379 557 -373
rect 691 -379 749 -373
<< pwell >>
rect -995 441 995 475
rect -995 -441 -961 441
rect 961 -441 995 441
rect -995 -475 995 -441
<< nmos >>
rect -831 109 -801 301
rect -735 109 -705 301
rect -639 109 -609 301
rect -543 109 -513 301
rect -447 109 -417 301
rect -351 109 -321 301
rect -255 109 -225 301
rect -159 109 -129 301
rect -63 109 -33 301
rect 33 109 63 301
rect 129 109 159 301
rect 225 109 255 301
rect 321 109 351 301
rect 417 109 447 301
rect 513 109 543 301
rect 609 109 639 301
rect 705 109 735 301
rect 801 109 831 301
rect -831 -301 -801 -109
rect -735 -301 -705 -109
rect -639 -301 -609 -109
rect -543 -301 -513 -109
rect -447 -301 -417 -109
rect -351 -301 -321 -109
rect -255 -301 -225 -109
rect -159 -301 -129 -109
rect -63 -301 -33 -109
rect 33 -301 63 -109
rect 129 -301 159 -109
rect 225 -301 255 -109
rect 321 -301 351 -109
rect 417 -301 447 -109
rect 513 -301 543 -109
rect 609 -301 639 -109
rect 705 -301 735 -109
rect 801 -301 831 -109
<< ndiff >>
rect -893 256 -831 301
rect -893 222 -881 256
rect -847 222 -831 256
rect -893 188 -831 222
rect -893 154 -881 188
rect -847 154 -831 188
rect -893 109 -831 154
rect -801 256 -735 301
rect -801 222 -785 256
rect -751 222 -735 256
rect -801 188 -735 222
rect -801 154 -785 188
rect -751 154 -735 188
rect -801 109 -735 154
rect -705 256 -639 301
rect -705 222 -689 256
rect -655 222 -639 256
rect -705 188 -639 222
rect -705 154 -689 188
rect -655 154 -639 188
rect -705 109 -639 154
rect -609 256 -543 301
rect -609 222 -593 256
rect -559 222 -543 256
rect -609 188 -543 222
rect -609 154 -593 188
rect -559 154 -543 188
rect -609 109 -543 154
rect -513 256 -447 301
rect -513 222 -497 256
rect -463 222 -447 256
rect -513 188 -447 222
rect -513 154 -497 188
rect -463 154 -447 188
rect -513 109 -447 154
rect -417 256 -351 301
rect -417 222 -401 256
rect -367 222 -351 256
rect -417 188 -351 222
rect -417 154 -401 188
rect -367 154 -351 188
rect -417 109 -351 154
rect -321 256 -255 301
rect -321 222 -305 256
rect -271 222 -255 256
rect -321 188 -255 222
rect -321 154 -305 188
rect -271 154 -255 188
rect -321 109 -255 154
rect -225 256 -159 301
rect -225 222 -209 256
rect -175 222 -159 256
rect -225 188 -159 222
rect -225 154 -209 188
rect -175 154 -159 188
rect -225 109 -159 154
rect -129 256 -63 301
rect -129 222 -113 256
rect -79 222 -63 256
rect -129 188 -63 222
rect -129 154 -113 188
rect -79 154 -63 188
rect -129 109 -63 154
rect -33 256 33 301
rect -33 222 -17 256
rect 17 222 33 256
rect -33 188 33 222
rect -33 154 -17 188
rect 17 154 33 188
rect -33 109 33 154
rect 63 256 129 301
rect 63 222 79 256
rect 113 222 129 256
rect 63 188 129 222
rect 63 154 79 188
rect 113 154 129 188
rect 63 109 129 154
rect 159 256 225 301
rect 159 222 175 256
rect 209 222 225 256
rect 159 188 225 222
rect 159 154 175 188
rect 209 154 225 188
rect 159 109 225 154
rect 255 256 321 301
rect 255 222 271 256
rect 305 222 321 256
rect 255 188 321 222
rect 255 154 271 188
rect 305 154 321 188
rect 255 109 321 154
rect 351 256 417 301
rect 351 222 367 256
rect 401 222 417 256
rect 351 188 417 222
rect 351 154 367 188
rect 401 154 417 188
rect 351 109 417 154
rect 447 256 513 301
rect 447 222 463 256
rect 497 222 513 256
rect 447 188 513 222
rect 447 154 463 188
rect 497 154 513 188
rect 447 109 513 154
rect 543 256 609 301
rect 543 222 559 256
rect 593 222 609 256
rect 543 188 609 222
rect 543 154 559 188
rect 593 154 609 188
rect 543 109 609 154
rect 639 256 705 301
rect 639 222 655 256
rect 689 222 705 256
rect 639 188 705 222
rect 639 154 655 188
rect 689 154 705 188
rect 639 109 705 154
rect 735 256 801 301
rect 735 222 751 256
rect 785 222 801 256
rect 735 188 801 222
rect 735 154 751 188
rect 785 154 801 188
rect 735 109 801 154
rect 831 256 893 301
rect 831 222 847 256
rect 881 222 893 256
rect 831 188 893 222
rect 831 154 847 188
rect 881 154 893 188
rect 831 109 893 154
rect -893 -154 -831 -109
rect -893 -188 -881 -154
rect -847 -188 -831 -154
rect -893 -222 -831 -188
rect -893 -256 -881 -222
rect -847 -256 -831 -222
rect -893 -301 -831 -256
rect -801 -154 -735 -109
rect -801 -188 -785 -154
rect -751 -188 -735 -154
rect -801 -222 -735 -188
rect -801 -256 -785 -222
rect -751 -256 -735 -222
rect -801 -301 -735 -256
rect -705 -154 -639 -109
rect -705 -188 -689 -154
rect -655 -188 -639 -154
rect -705 -222 -639 -188
rect -705 -256 -689 -222
rect -655 -256 -639 -222
rect -705 -301 -639 -256
rect -609 -154 -543 -109
rect -609 -188 -593 -154
rect -559 -188 -543 -154
rect -609 -222 -543 -188
rect -609 -256 -593 -222
rect -559 -256 -543 -222
rect -609 -301 -543 -256
rect -513 -154 -447 -109
rect -513 -188 -497 -154
rect -463 -188 -447 -154
rect -513 -222 -447 -188
rect -513 -256 -497 -222
rect -463 -256 -447 -222
rect -513 -301 -447 -256
rect -417 -154 -351 -109
rect -417 -188 -401 -154
rect -367 -188 -351 -154
rect -417 -222 -351 -188
rect -417 -256 -401 -222
rect -367 -256 -351 -222
rect -417 -301 -351 -256
rect -321 -154 -255 -109
rect -321 -188 -305 -154
rect -271 -188 -255 -154
rect -321 -222 -255 -188
rect -321 -256 -305 -222
rect -271 -256 -255 -222
rect -321 -301 -255 -256
rect -225 -154 -159 -109
rect -225 -188 -209 -154
rect -175 -188 -159 -154
rect -225 -222 -159 -188
rect -225 -256 -209 -222
rect -175 -256 -159 -222
rect -225 -301 -159 -256
rect -129 -154 -63 -109
rect -129 -188 -113 -154
rect -79 -188 -63 -154
rect -129 -222 -63 -188
rect -129 -256 -113 -222
rect -79 -256 -63 -222
rect -129 -301 -63 -256
rect -33 -154 33 -109
rect -33 -188 -17 -154
rect 17 -188 33 -154
rect -33 -222 33 -188
rect -33 -256 -17 -222
rect 17 -256 33 -222
rect -33 -301 33 -256
rect 63 -154 129 -109
rect 63 -188 79 -154
rect 113 -188 129 -154
rect 63 -222 129 -188
rect 63 -256 79 -222
rect 113 -256 129 -222
rect 63 -301 129 -256
rect 159 -154 225 -109
rect 159 -188 175 -154
rect 209 -188 225 -154
rect 159 -222 225 -188
rect 159 -256 175 -222
rect 209 -256 225 -222
rect 159 -301 225 -256
rect 255 -154 321 -109
rect 255 -188 271 -154
rect 305 -188 321 -154
rect 255 -222 321 -188
rect 255 -256 271 -222
rect 305 -256 321 -222
rect 255 -301 321 -256
rect 351 -154 417 -109
rect 351 -188 367 -154
rect 401 -188 417 -154
rect 351 -222 417 -188
rect 351 -256 367 -222
rect 401 -256 417 -222
rect 351 -301 417 -256
rect 447 -154 513 -109
rect 447 -188 463 -154
rect 497 -188 513 -154
rect 447 -222 513 -188
rect 447 -256 463 -222
rect 497 -256 513 -222
rect 447 -301 513 -256
rect 543 -154 609 -109
rect 543 -188 559 -154
rect 593 -188 609 -154
rect 543 -222 609 -188
rect 543 -256 559 -222
rect 593 -256 609 -222
rect 543 -301 609 -256
rect 639 -154 705 -109
rect 639 -188 655 -154
rect 689 -188 705 -154
rect 639 -222 705 -188
rect 639 -256 655 -222
rect 689 -256 705 -222
rect 639 -301 705 -256
rect 735 -154 801 -109
rect 735 -188 751 -154
rect 785 -188 801 -154
rect 735 -222 801 -188
rect 735 -256 751 -222
rect 785 -256 801 -222
rect 735 -301 801 -256
rect 831 -154 893 -109
rect 831 -188 847 -154
rect 881 -188 893 -154
rect 831 -222 893 -188
rect 831 -256 847 -222
rect 881 -256 893 -222
rect 831 -301 893 -256
<< ndiffc >>
rect -881 222 -847 256
rect -881 154 -847 188
rect -785 222 -751 256
rect -785 154 -751 188
rect -689 222 -655 256
rect -689 154 -655 188
rect -593 222 -559 256
rect -593 154 -559 188
rect -497 222 -463 256
rect -497 154 -463 188
rect -401 222 -367 256
rect -401 154 -367 188
rect -305 222 -271 256
rect -305 154 -271 188
rect -209 222 -175 256
rect -209 154 -175 188
rect -113 222 -79 256
rect -113 154 -79 188
rect -17 222 17 256
rect -17 154 17 188
rect 79 222 113 256
rect 79 154 113 188
rect 175 222 209 256
rect 175 154 209 188
rect 271 222 305 256
rect 271 154 305 188
rect 367 222 401 256
rect 367 154 401 188
rect 463 222 497 256
rect 463 154 497 188
rect 559 222 593 256
rect 559 154 593 188
rect 655 222 689 256
rect 655 154 689 188
rect 751 222 785 256
rect 751 154 785 188
rect 847 222 881 256
rect 847 154 881 188
rect -881 -188 -847 -154
rect -881 -256 -847 -222
rect -785 -188 -751 -154
rect -785 -256 -751 -222
rect -689 -188 -655 -154
rect -689 -256 -655 -222
rect -593 -188 -559 -154
rect -593 -256 -559 -222
rect -497 -188 -463 -154
rect -497 -256 -463 -222
rect -401 -188 -367 -154
rect -401 -256 -367 -222
rect -305 -188 -271 -154
rect -305 -256 -271 -222
rect -209 -188 -175 -154
rect -209 -256 -175 -222
rect -113 -188 -79 -154
rect -113 -256 -79 -222
rect -17 -188 17 -154
rect -17 -256 17 -222
rect 79 -188 113 -154
rect 79 -256 113 -222
rect 175 -188 209 -154
rect 175 -256 209 -222
rect 271 -188 305 -154
rect 271 -256 305 -222
rect 367 -188 401 -154
rect 367 -256 401 -222
rect 463 -188 497 -154
rect 463 -256 497 -222
rect 559 -188 593 -154
rect 559 -256 593 -222
rect 655 -188 689 -154
rect 655 -256 689 -222
rect 751 -188 785 -154
rect 751 -256 785 -222
rect 847 -188 881 -154
rect 847 -256 881 -222
<< psubdiff >>
rect -995 441 -867 475
rect -833 441 -799 475
rect -765 441 -731 475
rect -697 441 -663 475
rect -629 441 -595 475
rect -561 441 -527 475
rect -493 441 -459 475
rect -425 441 -391 475
rect -357 441 -323 475
rect -289 441 -255 475
rect -221 441 -187 475
rect -153 441 -119 475
rect -85 441 -51 475
rect -17 441 17 475
rect 51 441 85 475
rect 119 441 153 475
rect 187 441 221 475
rect 255 441 289 475
rect 323 441 357 475
rect 391 441 425 475
rect 459 441 493 475
rect 527 441 561 475
rect 595 441 629 475
rect 663 441 697 475
rect 731 441 765 475
rect 799 441 833 475
rect 867 441 995 475
rect -995 357 -961 441
rect -995 289 -961 323
rect 961 357 995 441
rect -995 221 -961 255
rect -995 153 -961 187
rect -995 85 -961 119
rect 961 289 995 323
rect 961 221 995 255
rect 961 153 995 187
rect -995 17 -961 51
rect 961 85 995 119
rect -995 -51 -961 -17
rect 961 17 995 51
rect -995 -119 -961 -85
rect 961 -51 995 -17
rect -995 -187 -961 -153
rect -995 -255 -961 -221
rect -995 -323 -961 -289
rect 961 -119 995 -85
rect 961 -187 995 -153
rect 961 -255 995 -221
rect -995 -441 -961 -357
rect 961 -323 995 -289
rect 961 -441 995 -357
rect -995 -475 -867 -441
rect -833 -475 -799 -441
rect -765 -475 -731 -441
rect -697 -475 -663 -441
rect -629 -475 -595 -441
rect -561 -475 -527 -441
rect -493 -475 -459 -441
rect -425 -475 -391 -441
rect -357 -475 -323 -441
rect -289 -475 -255 -441
rect -221 -475 -187 -441
rect -153 -475 -119 -441
rect -85 -475 -51 -441
rect -17 -475 17 -441
rect 51 -475 85 -441
rect 119 -475 153 -441
rect 187 -475 221 -441
rect 255 -475 289 -441
rect 323 -475 357 -441
rect 391 -475 425 -441
rect 459 -475 493 -441
rect 527 -475 561 -441
rect 595 -475 629 -441
rect 663 -475 697 -441
rect 731 -475 765 -441
rect 799 -475 833 -441
rect 867 -475 995 -441
<< psubdiffcont >>
rect -867 441 -833 475
rect -799 441 -765 475
rect -731 441 -697 475
rect -663 441 -629 475
rect -595 441 -561 475
rect -527 441 -493 475
rect -459 441 -425 475
rect -391 441 -357 475
rect -323 441 -289 475
rect -255 441 -221 475
rect -187 441 -153 475
rect -119 441 -85 475
rect -51 441 -17 475
rect 17 441 51 475
rect 85 441 119 475
rect 153 441 187 475
rect 221 441 255 475
rect 289 441 323 475
rect 357 441 391 475
rect 425 441 459 475
rect 493 441 527 475
rect 561 441 595 475
rect 629 441 663 475
rect 697 441 731 475
rect 765 441 799 475
rect 833 441 867 475
rect -995 323 -961 357
rect 961 323 995 357
rect -995 255 -961 289
rect -995 187 -961 221
rect -995 119 -961 153
rect 961 255 995 289
rect 961 187 995 221
rect 961 119 995 153
rect -995 51 -961 85
rect 961 51 995 85
rect -995 -17 -961 17
rect 961 -17 995 17
rect -995 -85 -961 -51
rect 961 -85 995 -51
rect -995 -153 -961 -119
rect -995 -221 -961 -187
rect -995 -289 -961 -255
rect 961 -153 995 -119
rect 961 -221 995 -187
rect 961 -289 995 -255
rect -995 -357 -961 -323
rect 961 -357 995 -323
rect -867 -475 -833 -441
rect -799 -475 -765 -441
rect -731 -475 -697 -441
rect -663 -475 -629 -441
rect -595 -475 -561 -441
rect -527 -475 -493 -441
rect -459 -475 -425 -441
rect -391 -475 -357 -441
rect -323 -475 -289 -441
rect -255 -475 -221 -441
rect -187 -475 -153 -441
rect -119 -475 -85 -441
rect -51 -475 -17 -441
rect 17 -475 51 -441
rect 85 -475 119 -441
rect 153 -475 187 -441
rect 221 -475 255 -441
rect 289 -475 323 -441
rect 357 -475 391 -441
rect 425 -475 459 -441
rect 493 -475 527 -441
rect 561 -475 595 -441
rect 629 -475 663 -441
rect 697 -475 731 -441
rect 765 -475 799 -441
rect 833 -475 867 -441
<< poly >>
rect -849 373 -783 389
rect -849 339 -833 373
rect -799 339 -783 373
rect -849 323 -783 339
rect -657 373 -591 389
rect -657 339 -641 373
rect -607 339 -591 373
rect -831 301 -801 323
rect -735 301 -705 327
rect -657 323 -591 339
rect -465 373 -399 389
rect -465 339 -449 373
rect -415 339 -399 373
rect -639 301 -609 323
rect -543 301 -513 327
rect -465 323 -399 339
rect -273 373 -207 389
rect -273 339 -257 373
rect -223 339 -207 373
rect -447 301 -417 323
rect -351 301 -321 327
rect -273 323 -207 339
rect -81 373 -15 389
rect -81 339 -65 373
rect -31 339 -15 373
rect -255 301 -225 323
rect -159 301 -129 327
rect -81 323 -15 339
rect 111 373 177 389
rect 111 339 127 373
rect 161 339 177 373
rect -63 301 -33 323
rect 33 301 63 327
rect 111 323 177 339
rect 303 373 369 389
rect 303 339 319 373
rect 353 339 369 373
rect 129 301 159 323
rect 225 301 255 327
rect 303 323 369 339
rect 495 373 561 389
rect 495 339 511 373
rect 545 339 561 373
rect 321 301 351 323
rect 417 301 447 327
rect 495 323 561 339
rect 687 373 753 389
rect 687 339 703 373
rect 737 339 753 373
rect 513 301 543 323
rect 609 301 639 327
rect 687 323 753 339
rect 705 301 735 323
rect 801 301 831 327
rect -831 83 -801 109
rect -735 87 -705 109
rect -753 71 -687 87
rect -639 83 -609 109
rect -543 87 -513 109
rect -753 37 -737 71
rect -703 37 -687 71
rect -753 21 -687 37
rect -561 71 -495 87
rect -447 83 -417 109
rect -351 87 -321 109
rect -561 37 -545 71
rect -511 37 -495 71
rect -561 21 -495 37
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 513 83 543 109
rect 609 87 639 109
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect 591 71 657 87
rect 705 83 735 109
rect 801 87 831 109
rect 591 37 607 71
rect 641 37 657 71
rect 591 21 657 37
rect 783 71 849 87
rect 783 37 799 71
rect 833 37 849 71
rect 783 21 849 37
rect -753 -37 -687 -21
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -831 -109 -801 -83
rect -753 -87 -687 -71
rect -561 -37 -495 -21
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -735 -109 -705 -87
rect -639 -109 -609 -83
rect -561 -87 -495 -71
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -543 -109 -513 -87
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 591 -37 657 -21
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 417 -109 447 -87
rect 513 -109 543 -83
rect 591 -87 657 -71
rect 783 -37 849 -21
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 609 -109 639 -87
rect 705 -109 735 -83
rect 783 -87 849 -71
rect 801 -109 831 -87
rect -831 -323 -801 -301
rect -849 -339 -783 -323
rect -735 -327 -705 -301
rect -639 -323 -609 -301
rect -849 -373 -833 -339
rect -799 -373 -783 -339
rect -849 -389 -783 -373
rect -657 -339 -591 -323
rect -543 -327 -513 -301
rect -447 -323 -417 -301
rect -657 -373 -641 -339
rect -607 -373 -591 -339
rect -657 -389 -591 -373
rect -465 -339 -399 -323
rect -351 -327 -321 -301
rect -255 -323 -225 -301
rect -465 -373 -449 -339
rect -415 -373 -399 -339
rect -465 -389 -399 -373
rect -273 -339 -207 -323
rect -159 -327 -129 -301
rect -63 -323 -33 -301
rect -273 -373 -257 -339
rect -223 -373 -207 -339
rect -273 -389 -207 -373
rect -81 -339 -15 -323
rect 33 -327 63 -301
rect 129 -323 159 -301
rect -81 -373 -65 -339
rect -31 -373 -15 -339
rect -81 -389 -15 -373
rect 111 -339 177 -323
rect 225 -327 255 -301
rect 321 -323 351 -301
rect 111 -373 127 -339
rect 161 -373 177 -339
rect 111 -389 177 -373
rect 303 -339 369 -323
rect 417 -327 447 -301
rect 513 -323 543 -301
rect 303 -373 319 -339
rect 353 -373 369 -339
rect 303 -389 369 -373
rect 495 -339 561 -323
rect 609 -327 639 -301
rect 705 -323 735 -301
rect 495 -373 511 -339
rect 545 -373 561 -339
rect 495 -389 561 -373
rect 687 -339 753 -323
rect 801 -327 831 -301
rect 687 -373 703 -339
rect 737 -373 753 -339
rect 687 -389 753 -373
<< polycont >>
rect -833 339 -799 373
rect -641 339 -607 373
rect -449 339 -415 373
rect -257 339 -223 373
rect -65 339 -31 373
rect 127 339 161 373
rect 319 339 353 373
rect 511 339 545 373
rect 703 339 737 373
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect -833 -373 -799 -339
rect -641 -373 -607 -339
rect -449 -373 -415 -339
rect -257 -373 -223 -339
rect -65 -373 -31 -339
rect 127 -373 161 -339
rect 319 -373 353 -339
rect 511 -373 545 -339
rect 703 -373 737 -339
<< locali >>
rect -995 441 -867 475
rect -833 441 -799 475
rect -765 441 -731 475
rect -697 441 -663 475
rect -629 441 -595 475
rect -561 441 -527 475
rect -493 441 -459 475
rect -425 441 -391 475
rect -357 441 -323 475
rect -289 441 -255 475
rect -221 441 -187 475
rect -153 441 -119 475
rect -85 441 -51 475
rect -17 441 17 475
rect 51 441 85 475
rect 119 441 153 475
rect 187 441 221 475
rect 255 441 289 475
rect 323 441 357 475
rect 391 441 425 475
rect 459 441 493 475
rect 527 441 561 475
rect 595 441 629 475
rect 663 441 697 475
rect 731 441 765 475
rect 799 441 833 475
rect 867 441 995 475
rect -995 357 -961 441
rect -849 339 -833 373
rect -799 339 -783 373
rect -657 339 -641 373
rect -607 339 -591 373
rect -465 339 -449 373
rect -415 339 -399 373
rect -273 339 -257 373
rect -223 339 -207 373
rect -81 339 -65 373
rect -31 339 -15 373
rect 111 339 127 373
rect 161 339 177 373
rect 303 339 319 373
rect 353 339 369 373
rect 495 339 511 373
rect 545 339 561 373
rect 687 339 703 373
rect 737 339 753 373
rect 961 357 995 441
rect -995 289 -961 323
rect -995 221 -961 255
rect -995 153 -961 187
rect -995 85 -961 119
rect -881 258 -847 305
rect -881 188 -847 222
rect -881 105 -847 152
rect -785 258 -751 305
rect -785 188 -751 222
rect -785 105 -751 152
rect -689 258 -655 305
rect -689 188 -655 222
rect -689 105 -655 152
rect -593 258 -559 305
rect -593 188 -559 222
rect -593 105 -559 152
rect -497 258 -463 305
rect -497 188 -463 222
rect -497 105 -463 152
rect -401 258 -367 305
rect -401 188 -367 222
rect -401 105 -367 152
rect -305 258 -271 305
rect -305 188 -271 222
rect -305 105 -271 152
rect -209 258 -175 305
rect -209 188 -175 222
rect -209 105 -175 152
rect -113 258 -79 305
rect -113 188 -79 222
rect -113 105 -79 152
rect -17 258 17 305
rect -17 188 17 222
rect -17 105 17 152
rect 79 258 113 305
rect 79 188 113 222
rect 79 105 113 152
rect 175 258 209 305
rect 175 188 209 222
rect 175 105 209 152
rect 271 258 305 305
rect 271 188 305 222
rect 271 105 305 152
rect 367 258 401 305
rect 367 188 401 222
rect 367 105 401 152
rect 463 258 497 305
rect 463 188 497 222
rect 463 105 497 152
rect 559 258 593 305
rect 559 188 593 222
rect 559 105 593 152
rect 655 258 689 305
rect 655 188 689 222
rect 655 105 689 152
rect 751 258 785 305
rect 751 188 785 222
rect 751 105 785 152
rect 847 258 881 305
rect 847 188 881 222
rect 847 105 881 152
rect 961 289 995 323
rect 961 221 995 255
rect 961 153 995 187
rect 961 85 995 119
rect -995 17 -961 51
rect -753 37 -737 71
rect -703 37 -687 71
rect -561 37 -545 71
rect -511 37 -495 71
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect 591 37 607 71
rect 641 37 657 71
rect 783 37 799 71
rect 833 37 849 71
rect -995 -51 -961 -17
rect 961 17 995 51
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 961 -51 995 -17
rect -995 -119 -961 -85
rect -995 -187 -961 -153
rect -995 -255 -961 -221
rect -995 -323 -961 -289
rect -881 -152 -847 -105
rect -881 -222 -847 -188
rect -881 -305 -847 -258
rect -785 -152 -751 -105
rect -785 -222 -751 -188
rect -785 -305 -751 -258
rect -689 -152 -655 -105
rect -689 -222 -655 -188
rect -689 -305 -655 -258
rect -593 -152 -559 -105
rect -593 -222 -559 -188
rect -593 -305 -559 -258
rect -497 -152 -463 -105
rect -497 -222 -463 -188
rect -497 -305 -463 -258
rect -401 -152 -367 -105
rect -401 -222 -367 -188
rect -401 -305 -367 -258
rect -305 -152 -271 -105
rect -305 -222 -271 -188
rect -305 -305 -271 -258
rect -209 -152 -175 -105
rect -209 -222 -175 -188
rect -209 -305 -175 -258
rect -113 -152 -79 -105
rect -113 -222 -79 -188
rect -113 -305 -79 -258
rect -17 -152 17 -105
rect -17 -222 17 -188
rect -17 -305 17 -258
rect 79 -152 113 -105
rect 79 -222 113 -188
rect 79 -305 113 -258
rect 175 -152 209 -105
rect 175 -222 209 -188
rect 175 -305 209 -258
rect 271 -152 305 -105
rect 271 -222 305 -188
rect 271 -305 305 -258
rect 367 -152 401 -105
rect 367 -222 401 -188
rect 367 -305 401 -258
rect 463 -152 497 -105
rect 463 -222 497 -188
rect 463 -305 497 -258
rect 559 -152 593 -105
rect 559 -222 593 -188
rect 559 -305 593 -258
rect 655 -152 689 -105
rect 655 -222 689 -188
rect 655 -305 689 -258
rect 751 -152 785 -105
rect 751 -222 785 -188
rect 751 -305 785 -258
rect 847 -152 881 -105
rect 847 -222 881 -188
rect 847 -305 881 -258
rect 961 -119 995 -85
rect 961 -187 995 -153
rect 961 -255 995 -221
rect 961 -323 995 -289
rect -995 -441 -961 -357
rect -849 -373 -833 -339
rect -799 -373 -783 -339
rect -657 -373 -641 -339
rect -607 -373 -591 -339
rect -465 -373 -449 -339
rect -415 -373 -399 -339
rect -273 -373 -257 -339
rect -223 -373 -207 -339
rect -81 -373 -65 -339
rect -31 -373 -15 -339
rect 111 -373 127 -339
rect 161 -373 177 -339
rect 303 -373 319 -339
rect 353 -373 369 -339
rect 495 -373 511 -339
rect 545 -373 561 -339
rect 687 -373 703 -339
rect 737 -373 753 -339
rect 961 -441 995 -357
rect -995 -475 -867 -441
rect -833 -475 -799 -441
rect -765 -475 -731 -441
rect -697 -475 -663 -441
rect -629 -475 -595 -441
rect -561 -475 -527 -441
rect -493 -475 -459 -441
rect -425 -475 -391 -441
rect -357 -475 -323 -441
rect -289 -475 -255 -441
rect -221 -475 -187 -441
rect -153 -475 -119 -441
rect -85 -475 -51 -441
rect -17 -475 17 -441
rect 51 -475 85 -441
rect 119 -475 153 -441
rect 187 -475 221 -441
rect 255 -475 289 -441
rect 323 -475 357 -441
rect 391 -475 425 -441
rect 459 -475 493 -441
rect 527 -475 561 -441
rect 595 -475 629 -441
rect 663 -475 697 -441
rect 731 -475 765 -441
rect 799 -475 833 -441
rect 867 -475 995 -441
<< viali >>
rect -833 339 -799 373
rect -641 339 -607 373
rect -449 339 -415 373
rect -257 339 -223 373
rect -65 339 -31 373
rect 127 339 161 373
rect 319 339 353 373
rect 511 339 545 373
rect 703 339 737 373
rect -881 256 -847 258
rect -881 224 -847 256
rect -881 154 -847 186
rect -881 152 -847 154
rect -785 256 -751 258
rect -785 224 -751 256
rect -785 154 -751 186
rect -785 152 -751 154
rect -689 256 -655 258
rect -689 224 -655 256
rect -689 154 -655 186
rect -689 152 -655 154
rect -593 256 -559 258
rect -593 224 -559 256
rect -593 154 -559 186
rect -593 152 -559 154
rect -497 256 -463 258
rect -497 224 -463 256
rect -497 154 -463 186
rect -497 152 -463 154
rect -401 256 -367 258
rect -401 224 -367 256
rect -401 154 -367 186
rect -401 152 -367 154
rect -305 256 -271 258
rect -305 224 -271 256
rect -305 154 -271 186
rect -305 152 -271 154
rect -209 256 -175 258
rect -209 224 -175 256
rect -209 154 -175 186
rect -209 152 -175 154
rect -113 256 -79 258
rect -113 224 -79 256
rect -113 154 -79 186
rect -113 152 -79 154
rect -17 256 17 258
rect -17 224 17 256
rect -17 154 17 186
rect -17 152 17 154
rect 79 256 113 258
rect 79 224 113 256
rect 79 154 113 186
rect 79 152 113 154
rect 175 256 209 258
rect 175 224 209 256
rect 175 154 209 186
rect 175 152 209 154
rect 271 256 305 258
rect 271 224 305 256
rect 271 154 305 186
rect 271 152 305 154
rect 367 256 401 258
rect 367 224 401 256
rect 367 154 401 186
rect 367 152 401 154
rect 463 256 497 258
rect 463 224 497 256
rect 463 154 497 186
rect 463 152 497 154
rect 559 256 593 258
rect 559 224 593 256
rect 559 154 593 186
rect 559 152 593 154
rect 655 256 689 258
rect 655 224 689 256
rect 655 154 689 186
rect 655 152 689 154
rect 751 256 785 258
rect 751 224 785 256
rect 751 154 785 186
rect 751 152 785 154
rect 847 256 881 258
rect 847 224 881 256
rect 847 154 881 186
rect 847 152 881 154
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect -881 -154 -847 -152
rect -881 -186 -847 -154
rect -881 -256 -847 -224
rect -881 -258 -847 -256
rect -785 -154 -751 -152
rect -785 -186 -751 -154
rect -785 -256 -751 -224
rect -785 -258 -751 -256
rect -689 -154 -655 -152
rect -689 -186 -655 -154
rect -689 -256 -655 -224
rect -689 -258 -655 -256
rect -593 -154 -559 -152
rect -593 -186 -559 -154
rect -593 -256 -559 -224
rect -593 -258 -559 -256
rect -497 -154 -463 -152
rect -497 -186 -463 -154
rect -497 -256 -463 -224
rect -497 -258 -463 -256
rect -401 -154 -367 -152
rect -401 -186 -367 -154
rect -401 -256 -367 -224
rect -401 -258 -367 -256
rect -305 -154 -271 -152
rect -305 -186 -271 -154
rect -305 -256 -271 -224
rect -305 -258 -271 -256
rect -209 -154 -175 -152
rect -209 -186 -175 -154
rect -209 -256 -175 -224
rect -209 -258 -175 -256
rect -113 -154 -79 -152
rect -113 -186 -79 -154
rect -113 -256 -79 -224
rect -113 -258 -79 -256
rect -17 -154 17 -152
rect -17 -186 17 -154
rect -17 -256 17 -224
rect -17 -258 17 -256
rect 79 -154 113 -152
rect 79 -186 113 -154
rect 79 -256 113 -224
rect 79 -258 113 -256
rect 175 -154 209 -152
rect 175 -186 209 -154
rect 175 -256 209 -224
rect 175 -258 209 -256
rect 271 -154 305 -152
rect 271 -186 305 -154
rect 271 -256 305 -224
rect 271 -258 305 -256
rect 367 -154 401 -152
rect 367 -186 401 -154
rect 367 -256 401 -224
rect 367 -258 401 -256
rect 463 -154 497 -152
rect 463 -186 497 -154
rect 463 -256 497 -224
rect 463 -258 497 -256
rect 559 -154 593 -152
rect 559 -186 593 -154
rect 559 -256 593 -224
rect 559 -258 593 -256
rect 655 -154 689 -152
rect 655 -186 689 -154
rect 655 -256 689 -224
rect 655 -258 689 -256
rect 751 -154 785 -152
rect 751 -186 785 -154
rect 751 -256 785 -224
rect 751 -258 785 -256
rect 847 -154 881 -152
rect 847 -186 881 -154
rect 847 -256 881 -224
rect 847 -258 881 -256
rect -833 -373 -799 -339
rect -641 -373 -607 -339
rect -449 -373 -415 -339
rect -257 -373 -223 -339
rect -65 -373 -31 -339
rect 127 -373 161 -339
rect 319 -373 353 -339
rect 511 -373 545 -339
rect 703 -373 737 -339
<< metal1 >>
rect -845 373 -787 379
rect -845 339 -833 373
rect -799 339 -787 373
rect -845 333 -787 339
rect -653 373 -595 379
rect -653 339 -641 373
rect -607 339 -595 373
rect -653 333 -595 339
rect -461 373 -403 379
rect -461 339 -449 373
rect -415 339 -403 373
rect -461 333 -403 339
rect -269 373 -211 379
rect -269 339 -257 373
rect -223 339 -211 373
rect -269 333 -211 339
rect -77 373 -19 379
rect -77 339 -65 373
rect -31 339 -19 373
rect -77 333 -19 339
rect 115 373 173 379
rect 115 339 127 373
rect 161 339 173 373
rect 115 333 173 339
rect 307 373 365 379
rect 307 339 319 373
rect 353 339 365 373
rect 307 333 365 339
rect 499 373 557 379
rect 499 339 511 373
rect 545 339 557 373
rect 499 333 557 339
rect 691 373 749 379
rect 691 339 703 373
rect 737 339 749 373
rect 691 333 749 339
rect -887 258 -841 301
rect -887 224 -881 258
rect -847 224 -841 258
rect -887 186 -841 224
rect -887 152 -881 186
rect -847 152 -841 186
rect -887 109 -841 152
rect -791 258 -745 301
rect -791 224 -785 258
rect -751 224 -745 258
rect -791 186 -745 224
rect -791 152 -785 186
rect -751 152 -745 186
rect -791 109 -745 152
rect -695 258 -649 301
rect -695 224 -689 258
rect -655 224 -649 258
rect -695 186 -649 224
rect -695 152 -689 186
rect -655 152 -649 186
rect -695 109 -649 152
rect -599 258 -553 301
rect -599 224 -593 258
rect -559 224 -553 258
rect -599 186 -553 224
rect -599 152 -593 186
rect -559 152 -553 186
rect -599 109 -553 152
rect -503 258 -457 301
rect -503 224 -497 258
rect -463 224 -457 258
rect -503 186 -457 224
rect -503 152 -497 186
rect -463 152 -457 186
rect -503 109 -457 152
rect -407 258 -361 301
rect -407 224 -401 258
rect -367 224 -361 258
rect -407 186 -361 224
rect -407 152 -401 186
rect -367 152 -361 186
rect -407 109 -361 152
rect -311 258 -265 301
rect -311 224 -305 258
rect -271 224 -265 258
rect -311 186 -265 224
rect -311 152 -305 186
rect -271 152 -265 186
rect -311 109 -265 152
rect -215 258 -169 301
rect -215 224 -209 258
rect -175 224 -169 258
rect -215 186 -169 224
rect -215 152 -209 186
rect -175 152 -169 186
rect -215 109 -169 152
rect -119 258 -73 301
rect -119 224 -113 258
rect -79 224 -73 258
rect -119 186 -73 224
rect -119 152 -113 186
rect -79 152 -73 186
rect -119 109 -73 152
rect -23 258 23 301
rect -23 224 -17 258
rect 17 224 23 258
rect -23 186 23 224
rect -23 152 -17 186
rect 17 152 23 186
rect -23 109 23 152
rect 73 258 119 301
rect 73 224 79 258
rect 113 224 119 258
rect 73 186 119 224
rect 73 152 79 186
rect 113 152 119 186
rect 73 109 119 152
rect 169 258 215 301
rect 169 224 175 258
rect 209 224 215 258
rect 169 186 215 224
rect 169 152 175 186
rect 209 152 215 186
rect 169 109 215 152
rect 265 258 311 301
rect 265 224 271 258
rect 305 224 311 258
rect 265 186 311 224
rect 265 152 271 186
rect 305 152 311 186
rect 265 109 311 152
rect 361 258 407 301
rect 361 224 367 258
rect 401 224 407 258
rect 361 186 407 224
rect 361 152 367 186
rect 401 152 407 186
rect 361 109 407 152
rect 457 258 503 301
rect 457 224 463 258
rect 497 224 503 258
rect 457 186 503 224
rect 457 152 463 186
rect 497 152 503 186
rect 457 109 503 152
rect 553 258 599 301
rect 553 224 559 258
rect 593 224 599 258
rect 553 186 599 224
rect 553 152 559 186
rect 593 152 599 186
rect 553 109 599 152
rect 649 258 695 301
rect 649 224 655 258
rect 689 224 695 258
rect 649 186 695 224
rect 649 152 655 186
rect 689 152 695 186
rect 649 109 695 152
rect 745 258 791 301
rect 745 224 751 258
rect 785 224 791 258
rect 745 186 791 224
rect 745 152 751 186
rect 785 152 791 186
rect 745 109 791 152
rect 841 258 887 301
rect 841 224 847 258
rect 881 224 887 258
rect 841 186 887 224
rect 841 152 847 186
rect 881 152 887 186
rect 841 109 887 152
rect -749 71 -691 77
rect -749 37 -737 71
rect -703 37 -691 71
rect -749 31 -691 37
rect -557 71 -499 77
rect -557 37 -545 71
rect -511 37 -499 71
rect -557 31 -499 37
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect 595 71 653 77
rect 595 37 607 71
rect 641 37 653 71
rect 595 31 653 37
rect 787 71 845 77
rect 787 37 799 71
rect 833 37 845 71
rect 787 31 845 37
rect -749 -37 -691 -31
rect -749 -71 -737 -37
rect -703 -71 -691 -37
rect -749 -77 -691 -71
rect -557 -37 -499 -31
rect -557 -71 -545 -37
rect -511 -71 -499 -37
rect -557 -77 -499 -71
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect 595 -37 653 -31
rect 595 -71 607 -37
rect 641 -71 653 -37
rect 595 -77 653 -71
rect 787 -37 845 -31
rect 787 -71 799 -37
rect 833 -71 845 -37
rect 787 -77 845 -71
rect -887 -152 -841 -109
rect -887 -186 -881 -152
rect -847 -186 -841 -152
rect -887 -224 -841 -186
rect -887 -258 -881 -224
rect -847 -258 -841 -224
rect -887 -301 -841 -258
rect -791 -152 -745 -109
rect -791 -186 -785 -152
rect -751 -186 -745 -152
rect -791 -224 -745 -186
rect -791 -258 -785 -224
rect -751 -258 -745 -224
rect -791 -301 -745 -258
rect -695 -152 -649 -109
rect -695 -186 -689 -152
rect -655 -186 -649 -152
rect -695 -224 -649 -186
rect -695 -258 -689 -224
rect -655 -258 -649 -224
rect -695 -301 -649 -258
rect -599 -152 -553 -109
rect -599 -186 -593 -152
rect -559 -186 -553 -152
rect -599 -224 -553 -186
rect -599 -258 -593 -224
rect -559 -258 -553 -224
rect -599 -301 -553 -258
rect -503 -152 -457 -109
rect -503 -186 -497 -152
rect -463 -186 -457 -152
rect -503 -224 -457 -186
rect -503 -258 -497 -224
rect -463 -258 -457 -224
rect -503 -301 -457 -258
rect -407 -152 -361 -109
rect -407 -186 -401 -152
rect -367 -186 -361 -152
rect -407 -224 -361 -186
rect -407 -258 -401 -224
rect -367 -258 -361 -224
rect -407 -301 -361 -258
rect -311 -152 -265 -109
rect -311 -186 -305 -152
rect -271 -186 -265 -152
rect -311 -224 -265 -186
rect -311 -258 -305 -224
rect -271 -258 -265 -224
rect -311 -301 -265 -258
rect -215 -152 -169 -109
rect -215 -186 -209 -152
rect -175 -186 -169 -152
rect -215 -224 -169 -186
rect -215 -258 -209 -224
rect -175 -258 -169 -224
rect -215 -301 -169 -258
rect -119 -152 -73 -109
rect -119 -186 -113 -152
rect -79 -186 -73 -152
rect -119 -224 -73 -186
rect -119 -258 -113 -224
rect -79 -258 -73 -224
rect -119 -301 -73 -258
rect -23 -152 23 -109
rect -23 -186 -17 -152
rect 17 -186 23 -152
rect -23 -224 23 -186
rect -23 -258 -17 -224
rect 17 -258 23 -224
rect -23 -301 23 -258
rect 73 -152 119 -109
rect 73 -186 79 -152
rect 113 -186 119 -152
rect 73 -224 119 -186
rect 73 -258 79 -224
rect 113 -258 119 -224
rect 73 -301 119 -258
rect 169 -152 215 -109
rect 169 -186 175 -152
rect 209 -186 215 -152
rect 169 -224 215 -186
rect 169 -258 175 -224
rect 209 -258 215 -224
rect 169 -301 215 -258
rect 265 -152 311 -109
rect 265 -186 271 -152
rect 305 -186 311 -152
rect 265 -224 311 -186
rect 265 -258 271 -224
rect 305 -258 311 -224
rect 265 -301 311 -258
rect 361 -152 407 -109
rect 361 -186 367 -152
rect 401 -186 407 -152
rect 361 -224 407 -186
rect 361 -258 367 -224
rect 401 -258 407 -224
rect 361 -301 407 -258
rect 457 -152 503 -109
rect 457 -186 463 -152
rect 497 -186 503 -152
rect 457 -224 503 -186
rect 457 -258 463 -224
rect 497 -258 503 -224
rect 457 -301 503 -258
rect 553 -152 599 -109
rect 553 -186 559 -152
rect 593 -186 599 -152
rect 553 -224 599 -186
rect 553 -258 559 -224
rect 593 -258 599 -224
rect 553 -301 599 -258
rect 649 -152 695 -109
rect 649 -186 655 -152
rect 689 -186 695 -152
rect 649 -224 695 -186
rect 649 -258 655 -224
rect 689 -258 695 -224
rect 649 -301 695 -258
rect 745 -152 791 -109
rect 745 -186 751 -152
rect 785 -186 791 -152
rect 745 -224 791 -186
rect 745 -258 751 -224
rect 785 -258 791 -224
rect 745 -301 791 -258
rect 841 -152 887 -109
rect 841 -186 847 -152
rect 881 -186 887 -152
rect 841 -224 887 -186
rect 841 -258 847 -224
rect 881 -258 887 -224
rect 841 -301 887 -258
rect -845 -339 -787 -333
rect -845 -373 -833 -339
rect -799 -373 -787 -339
rect -845 -379 -787 -373
rect -653 -339 -595 -333
rect -653 -373 -641 -339
rect -607 -373 -595 -339
rect -653 -379 -595 -373
rect -461 -339 -403 -333
rect -461 -373 -449 -339
rect -415 -373 -403 -339
rect -461 -379 -403 -373
rect -269 -339 -211 -333
rect -269 -373 -257 -339
rect -223 -373 -211 -339
rect -269 -379 -211 -373
rect -77 -339 -19 -333
rect -77 -373 -65 -339
rect -31 -373 -19 -339
rect -77 -379 -19 -373
rect 115 -339 173 -333
rect 115 -373 127 -339
rect 161 -373 173 -339
rect 115 -379 173 -373
rect 307 -339 365 -333
rect 307 -373 319 -339
rect 353 -373 365 -339
rect 307 -379 365 -373
rect 499 -339 557 -333
rect 499 -373 511 -339
rect 545 -373 557 -339
rect 499 -379 557 -373
rect 691 -339 749 -333
rect 691 -373 703 -339
rect 737 -373 749 -339
rect 691 -379 749 -373
<< properties >>
string FIXED_BBOX -978 -458 978 458
<< end >>
