magic
tech sky130A
magscale 1 2
timestamp 1627987662
<< nwell >>
rect 124 792 188 1230
rect 316 792 380 1230
rect 508 792 572 1230
rect 700 792 764 1230
rect 892 792 956 1230
rect 1084 792 1148 1230
rect 1276 792 1340 1230
rect 1468 792 1532 1230
rect 1660 792 1724 1230
rect 124 114 188 552
rect 316 114 380 552
rect 508 114 572 552
rect 700 114 764 552
rect 892 114 956 552
rect 1084 114 1148 552
rect 1276 114 1340 552
rect 1468 114 1532 552
rect 1660 114 1724 552
<< pdiff >>
rect 124 1221 188 1230
rect 124 803 140 1221
rect 174 803 188 1221
rect 124 792 188 803
rect 316 1221 380 1230
rect 316 803 332 1221
rect 366 803 380 1221
rect 316 792 380 803
rect 508 1221 572 1230
rect 508 803 524 1221
rect 558 803 572 1221
rect 508 792 572 803
rect 700 1221 764 1230
rect 700 803 716 1221
rect 750 803 764 1221
rect 700 792 764 803
rect 892 1221 956 1230
rect 892 803 908 1221
rect 942 803 956 1221
rect 892 792 956 803
rect 1084 1221 1148 1230
rect 1084 803 1100 1221
rect 1134 803 1148 1221
rect 1084 792 1148 803
rect 1276 1221 1340 1230
rect 1276 803 1292 1221
rect 1326 803 1340 1221
rect 1276 792 1340 803
rect 1468 1221 1532 1230
rect 1468 803 1484 1221
rect 1518 803 1532 1221
rect 1468 792 1532 803
rect 1660 1221 1724 1230
rect 1660 803 1676 1221
rect 1710 803 1724 1221
rect 1660 792 1724 803
rect 124 543 188 552
rect 124 125 140 543
rect 174 125 188 543
rect 124 114 188 125
rect 316 543 380 552
rect 316 125 332 543
rect 366 125 380 543
rect 316 114 380 125
rect 508 543 572 552
rect 508 125 524 543
rect 558 125 572 543
rect 508 114 572 125
rect 700 543 764 552
rect 700 125 716 543
rect 750 125 764 543
rect 700 114 764 125
rect 892 543 956 552
rect 892 125 908 543
rect 942 125 956 543
rect 892 114 956 125
rect 1084 543 1148 552
rect 1084 125 1100 543
rect 1134 125 1148 543
rect 1084 114 1148 125
rect 1276 543 1340 552
rect 1276 125 1292 543
rect 1326 125 1340 543
rect 1276 114 1340 125
rect 1468 543 1532 552
rect 1468 125 1484 543
rect 1518 125 1532 543
rect 1468 114 1532 125
rect 1660 543 1724 552
rect 1660 125 1676 543
rect 1710 125 1724 543
rect 1660 114 1724 125
<< pdiffc >>
rect 140 803 174 1221
rect 332 803 366 1221
rect 524 803 558 1221
rect 716 803 750 1221
rect 908 803 942 1221
rect 1100 803 1134 1221
rect 1292 803 1326 1221
rect 1484 803 1518 1221
rect 1676 803 1710 1221
rect 140 125 174 543
rect 332 125 366 543
rect 524 125 558 543
rect 716 125 750 543
rect 908 125 942 543
rect 1100 125 1134 543
rect 1292 125 1326 543
rect 1484 125 1518 543
rect 1676 125 1710 543
<< poly >>
rect 1659 1289 1756 1315
rect 1665 1285 1756 1289
rect 1726 1233 1756 1285
rect 1726 59 1756 113
rect 1673 55 1756 59
rect 1663 29 1756 55
rect 1665 -305 1760 -279
rect 1675 -309 1760 -305
rect 1730 -340 1760 -309
rect 1730 -987 1760 -942
rect 1669 -1017 1760 -987
<< locali >>
rect -72 1536 1920 1538
rect -72 1474 -68 1536
rect 1912 1474 1920 1536
rect -72 1462 1920 1474
rect -70 1388 1920 1462
rect 140 1221 174 1230
rect 140 792 174 803
rect 332 1221 366 1230
rect 332 792 366 803
rect 524 1221 558 1230
rect 524 792 558 803
rect 716 1221 750 1230
rect 716 792 750 803
rect 908 1221 942 1230
rect 908 792 942 803
rect 1100 1221 1134 1230
rect 1100 792 1134 803
rect 1292 1221 1326 1230
rect 1292 792 1326 803
rect 1484 1221 1518 1230
rect 1484 792 1518 803
rect 1676 1221 1710 1230
rect 1676 792 1710 803
rect 140 543 174 552
rect 140 114 174 125
rect 332 543 366 552
rect 332 114 366 125
rect 524 543 558 552
rect 524 114 558 125
rect 716 543 750 552
rect 716 114 750 125
rect 908 543 942 552
rect 908 114 942 125
rect 1100 543 1134 552
rect 1100 114 1134 125
rect 1292 543 1326 552
rect 1292 114 1326 125
rect 1484 543 1518 552
rect 1484 114 1518 125
rect 1676 543 1710 552
rect 1676 114 1710 125
rect -74 -1158 1926 -1094
rect -66 -1166 1926 -1158
rect -66 -1200 -58 -1166
rect -64 -1230 -58 -1200
rect 1914 -1230 1926 -1166
rect -64 -1242 1926 -1230
<< viali >>
rect -68 1474 1912 1536
rect 140 803 174 1221
rect 332 803 366 1221
rect 524 803 558 1221
rect 716 803 750 1221
rect 908 803 942 1221
rect 1100 803 1134 1221
rect 1292 803 1326 1221
rect 1484 803 1518 1221
rect 1676 803 1710 1221
rect 140 125 174 543
rect 332 125 366 543
rect 524 125 558 543
rect 716 125 750 543
rect 908 125 942 543
rect 1100 125 1134 543
rect 1292 125 1326 543
rect 1484 125 1518 543
rect 1676 125 1710 543
rect -58 -1230 1914 -1166
<< metal1 >>
rect -84 1542 1924 1554
rect -84 1478 -76 1542
rect 1916 1478 1924 1542
rect -84 1474 -68 1478
rect 1912 1474 1924 1478
rect -84 1464 1924 1474
rect 78 1274 1676 1322
rect 30 1220 94 1226
rect 30 798 36 1220
rect 88 798 94 1220
rect 30 792 94 798
rect 124 1224 188 1230
rect 124 798 130 1224
rect 182 798 188 1224
rect 124 792 188 798
rect 222 1220 286 1226
rect 222 798 228 1220
rect 280 798 286 1220
rect 222 792 286 798
rect 316 1224 380 1230
rect 316 798 322 1224
rect 374 798 380 1224
rect 316 792 380 798
rect 414 1220 478 1226
rect 414 798 420 1220
rect 472 798 478 1220
rect 414 792 478 798
rect 508 1224 572 1230
rect 508 798 514 1224
rect 566 798 572 1224
rect 508 792 572 798
rect 606 1220 670 1226
rect 606 798 612 1220
rect 664 798 670 1220
rect 606 792 670 798
rect 700 1224 764 1230
rect 700 798 706 1224
rect 758 798 764 1224
rect 700 792 764 798
rect 798 1220 862 1226
rect 798 798 804 1220
rect 856 798 862 1220
rect 798 792 862 798
rect 892 1224 956 1230
rect 892 798 898 1224
rect 950 798 956 1224
rect 892 792 956 798
rect 990 1220 1054 1226
rect 990 798 996 1220
rect 1048 798 1054 1220
rect 990 792 1054 798
rect 1084 1224 1148 1230
rect 1084 798 1090 1224
rect 1142 798 1148 1224
rect 1084 792 1148 798
rect 1182 1220 1246 1226
rect 1182 798 1188 1220
rect 1240 798 1246 1220
rect 1182 792 1246 798
rect 1276 1224 1340 1230
rect 1276 798 1282 1224
rect 1334 798 1340 1224
rect 1276 792 1340 798
rect 1374 1220 1438 1226
rect 1374 798 1380 1220
rect 1432 798 1438 1220
rect 1374 792 1438 798
rect 1468 1224 1532 1230
rect 1468 798 1474 1224
rect 1526 798 1532 1224
rect 1468 792 1532 798
rect 1566 1220 1630 1226
rect 1566 798 1572 1220
rect 1624 798 1630 1220
rect 1566 792 1630 798
rect 1660 1224 1724 1230
rect 1660 798 1666 1224
rect 1718 798 1724 1224
rect 1660 792 1724 798
rect 1758 1220 1822 1226
rect 1758 798 1764 1220
rect 1816 798 1822 1220
rect 1758 792 1822 798
rect -166 596 1772 752
rect -166 -564 -10 596
rect 30 542 94 548
rect 30 120 36 542
rect 88 120 94 542
rect 30 114 94 120
rect 124 546 188 552
rect 124 120 130 546
rect 182 120 188 546
rect 124 114 188 120
rect 222 542 286 548
rect 222 120 228 542
rect 280 120 286 542
rect 222 114 286 120
rect 316 546 380 552
rect 316 120 322 546
rect 374 120 380 546
rect 316 114 380 120
rect 414 542 478 548
rect 414 120 420 542
rect 472 120 478 542
rect 414 114 478 120
rect 508 546 572 552
rect 508 120 514 546
rect 566 120 572 546
rect 508 114 572 120
rect 606 542 670 548
rect 606 120 612 542
rect 664 120 670 542
rect 606 114 670 120
rect 700 546 764 552
rect 700 120 706 546
rect 758 120 764 546
rect 700 114 764 120
rect 798 542 862 548
rect 798 120 804 542
rect 856 120 862 542
rect 798 114 862 120
rect 892 546 956 552
rect 892 120 898 546
rect 950 120 956 546
rect 892 114 956 120
rect 990 542 1054 548
rect 990 120 996 542
rect 1048 120 1054 542
rect 990 114 1054 120
rect 1084 546 1148 552
rect 1084 120 1090 546
rect 1142 120 1148 546
rect 1084 114 1148 120
rect 1182 542 1246 548
rect 1182 120 1188 542
rect 1240 120 1246 542
rect 1182 114 1246 120
rect 1276 546 1340 552
rect 1276 120 1282 546
rect 1334 120 1340 546
rect 1276 114 1340 120
rect 1374 542 1438 548
rect 1374 120 1380 542
rect 1432 120 1438 542
rect 1374 114 1438 120
rect 1468 546 1532 552
rect 1468 120 1474 546
rect 1526 120 1532 546
rect 1468 114 1532 120
rect 1566 542 1630 548
rect 1566 120 1572 542
rect 1624 120 1630 542
rect 1566 114 1630 120
rect 1660 546 1724 552
rect 1660 120 1666 546
rect 1718 120 1724 546
rect 1660 114 1724 120
rect 1758 542 1822 548
rect 1758 120 1764 542
rect 1816 120 1822 542
rect 1758 114 1822 120
rect 78 26 1676 74
rect 82 -308 1680 -260
rect 34 -350 98 -344
rect 34 -526 40 -350
rect 92 -526 98 -350
rect 34 -532 98 -526
rect 130 -350 194 -344
rect 130 -524 136 -350
rect 188 -524 194 -350
rect 130 -530 194 -524
rect 226 -350 290 -344
rect 226 -526 232 -350
rect 284 -526 290 -350
rect 226 -532 290 -526
rect 322 -350 386 -344
rect 322 -524 328 -350
rect 380 -524 386 -350
rect 322 -530 386 -524
rect 418 -350 482 -344
rect 418 -526 424 -350
rect 476 -526 482 -350
rect 418 -532 482 -526
rect 514 -350 578 -344
rect 514 -524 520 -350
rect 572 -524 578 -350
rect 514 -530 578 -524
rect 610 -350 674 -344
rect 610 -526 616 -350
rect 668 -526 674 -350
rect 610 -532 674 -526
rect 706 -350 770 -344
rect 706 -524 712 -350
rect 764 -524 770 -350
rect 706 -530 770 -524
rect 802 -350 866 -344
rect 802 -526 808 -350
rect 860 -526 866 -350
rect 802 -532 866 -526
rect 898 -350 962 -344
rect 898 -524 904 -350
rect 956 -524 962 -350
rect 898 -530 962 -524
rect 994 -350 1058 -344
rect 994 -526 1000 -350
rect 1052 -526 1058 -350
rect 994 -532 1058 -526
rect 1090 -350 1154 -344
rect 1090 -524 1096 -350
rect 1148 -524 1154 -350
rect 1090 -530 1154 -524
rect 1186 -350 1250 -344
rect 1186 -526 1192 -350
rect 1244 -526 1250 -350
rect 1186 -532 1250 -526
rect 1282 -350 1346 -344
rect 1282 -524 1288 -350
rect 1340 -524 1346 -350
rect 1282 -530 1346 -524
rect 1378 -350 1442 -344
rect 1378 -526 1384 -350
rect 1436 -526 1442 -350
rect 1378 -532 1442 -526
rect 1474 -350 1538 -344
rect 1474 -524 1480 -350
rect 1532 -524 1538 -350
rect 1474 -530 1538 -524
rect 1570 -350 1634 -344
rect 1570 -526 1576 -350
rect 1628 -526 1634 -350
rect 1570 -532 1634 -526
rect 1666 -350 1730 -344
rect 1666 -524 1672 -350
rect 1724 -524 1730 -350
rect 1666 -530 1730 -524
rect 1762 -350 1826 -344
rect 1762 -526 1768 -350
rect 1820 -526 1826 -350
rect 1762 -532 1826 -526
rect -166 -714 1776 -564
rect -163 -718 1776 -714
rect 34 -758 98 -752
rect 34 -934 40 -758
rect 92 -934 98 -758
rect 34 -940 98 -934
rect 130 -760 194 -754
rect 130 -934 136 -760
rect 188 -934 194 -760
rect 130 -940 194 -934
rect 226 -758 290 -752
rect 226 -934 232 -758
rect 284 -934 290 -758
rect 226 -940 290 -934
rect 322 -760 386 -754
rect 322 -934 328 -760
rect 380 -934 386 -760
rect 322 -940 386 -934
rect 418 -758 482 -752
rect 418 -934 424 -758
rect 476 -934 482 -758
rect 418 -940 482 -934
rect 514 -760 578 -754
rect 514 -934 520 -760
rect 572 -934 578 -760
rect 514 -940 578 -934
rect 610 -758 674 -752
rect 610 -934 616 -758
rect 668 -934 674 -758
rect 610 -940 674 -934
rect 706 -760 770 -754
rect 706 -934 712 -760
rect 764 -934 770 -760
rect 706 -940 770 -934
rect 802 -758 866 -752
rect 802 -934 808 -758
rect 860 -934 866 -758
rect 802 -940 866 -934
rect 898 -760 962 -754
rect 898 -934 904 -760
rect 956 -934 962 -760
rect 898 -940 962 -934
rect 994 -758 1058 -752
rect 994 -934 1000 -758
rect 1052 -934 1058 -758
rect 994 -940 1058 -934
rect 1090 -760 1154 -754
rect 1090 -934 1096 -760
rect 1148 -934 1154 -760
rect 1090 -940 1154 -934
rect 1186 -758 1250 -752
rect 1186 -934 1192 -758
rect 1244 -934 1250 -758
rect 1186 -940 1250 -934
rect 1282 -760 1346 -754
rect 1282 -934 1288 -760
rect 1340 -934 1346 -760
rect 1282 -940 1346 -934
rect 1378 -758 1442 -752
rect 1378 -934 1384 -758
rect 1436 -934 1442 -758
rect 1378 -940 1442 -934
rect 1474 -760 1538 -754
rect 1474 -934 1480 -760
rect 1532 -934 1538 -760
rect 1474 -940 1538 -934
rect 1570 -758 1634 -752
rect 1570 -934 1576 -758
rect 1628 -934 1634 -758
rect 1570 -940 1634 -934
rect 1666 -760 1730 -754
rect 1666 -934 1672 -760
rect 1724 -934 1730 -760
rect 1666 -940 1730 -934
rect 1762 -758 1826 -752
rect 1762 -934 1768 -758
rect 1820 -934 1826 -758
rect 1762 -940 1826 -934
rect 80 -1022 1730 -974
rect -76 -1148 1924 -1142
rect -76 -1150 1926 -1148
rect -76 -1234 -64 -1150
rect -74 -1238 -64 -1234
rect 1922 -1238 1926 -1150
rect -74 -1246 1926 -1238
<< via1 >>
rect -76 1536 1916 1542
rect -76 1478 -68 1536
rect -68 1478 1912 1536
rect 1912 1478 1916 1536
rect 36 798 88 1220
rect 130 1221 182 1224
rect 130 803 140 1221
rect 140 803 174 1221
rect 174 803 182 1221
rect 130 798 182 803
rect 228 798 280 1220
rect 322 1221 374 1224
rect 322 803 332 1221
rect 332 803 366 1221
rect 366 803 374 1221
rect 322 798 374 803
rect 420 798 472 1220
rect 514 1221 566 1224
rect 514 803 524 1221
rect 524 803 558 1221
rect 558 803 566 1221
rect 514 798 566 803
rect 612 798 664 1220
rect 706 1221 758 1224
rect 706 803 716 1221
rect 716 803 750 1221
rect 750 803 758 1221
rect 706 798 758 803
rect 804 798 856 1220
rect 898 1221 950 1224
rect 898 803 908 1221
rect 908 803 942 1221
rect 942 803 950 1221
rect 898 798 950 803
rect 996 798 1048 1220
rect 1090 1221 1142 1224
rect 1090 803 1100 1221
rect 1100 803 1134 1221
rect 1134 803 1142 1221
rect 1090 798 1142 803
rect 1188 798 1240 1220
rect 1282 1221 1334 1224
rect 1282 803 1292 1221
rect 1292 803 1326 1221
rect 1326 803 1334 1221
rect 1282 798 1334 803
rect 1380 798 1432 1220
rect 1474 1221 1526 1224
rect 1474 803 1484 1221
rect 1484 803 1518 1221
rect 1518 803 1526 1221
rect 1474 798 1526 803
rect 1572 798 1624 1220
rect 1666 1221 1718 1224
rect 1666 803 1676 1221
rect 1676 803 1710 1221
rect 1710 803 1718 1221
rect 1666 798 1718 803
rect 1764 798 1816 1220
rect 36 120 88 542
rect 130 543 182 546
rect 130 125 140 543
rect 140 125 174 543
rect 174 125 182 543
rect 130 120 182 125
rect 228 120 280 542
rect 322 543 374 546
rect 322 125 332 543
rect 332 125 366 543
rect 366 125 374 543
rect 322 120 374 125
rect 420 120 472 542
rect 514 543 566 546
rect 514 125 524 543
rect 524 125 558 543
rect 558 125 566 543
rect 514 120 566 125
rect 612 120 664 542
rect 706 543 758 546
rect 706 125 716 543
rect 716 125 750 543
rect 750 125 758 543
rect 706 120 758 125
rect 804 120 856 542
rect 898 543 950 546
rect 898 125 908 543
rect 908 125 942 543
rect 942 125 950 543
rect 898 120 950 125
rect 996 120 1048 542
rect 1090 543 1142 546
rect 1090 125 1100 543
rect 1100 125 1134 543
rect 1134 125 1142 543
rect 1090 120 1142 125
rect 1188 120 1240 542
rect 1282 543 1334 546
rect 1282 125 1292 543
rect 1292 125 1326 543
rect 1326 125 1334 543
rect 1282 120 1334 125
rect 1380 120 1432 542
rect 1474 543 1526 546
rect 1474 125 1484 543
rect 1484 125 1518 543
rect 1518 125 1526 543
rect 1474 120 1526 125
rect 1572 120 1624 542
rect 1666 543 1718 546
rect 1666 125 1676 543
rect 1676 125 1710 543
rect 1710 125 1718 543
rect 1666 120 1718 125
rect 1764 120 1816 542
rect 40 -526 92 -350
rect 136 -524 188 -350
rect 232 -526 284 -350
rect 328 -524 380 -350
rect 424 -526 476 -350
rect 520 -524 572 -350
rect 616 -526 668 -350
rect 712 -524 764 -350
rect 808 -526 860 -350
rect 904 -524 956 -350
rect 1000 -526 1052 -350
rect 1096 -524 1148 -350
rect 1192 -526 1244 -350
rect 1288 -524 1340 -350
rect 1384 -526 1436 -350
rect 1480 -524 1532 -350
rect 1576 -526 1628 -350
rect 1672 -524 1724 -350
rect 1768 -526 1820 -350
rect 40 -934 92 -758
rect 136 -934 188 -760
rect 232 -934 284 -758
rect 328 -934 380 -760
rect 424 -934 476 -758
rect 520 -934 572 -760
rect 616 -934 668 -758
rect 712 -934 764 -760
rect 808 -934 860 -758
rect 904 -934 956 -760
rect 1000 -934 1052 -758
rect 1096 -934 1148 -760
rect 1192 -934 1244 -758
rect 1288 -934 1340 -760
rect 1384 -934 1436 -758
rect 1480 -934 1532 -760
rect 1576 -934 1628 -758
rect 1672 -934 1724 -760
rect 1768 -934 1820 -758
rect -64 -1166 1922 -1150
rect -64 -1230 -58 -1166
rect -58 -1230 1914 -1166
rect 1914 -1230 1922 -1166
rect -64 -1238 1922 -1230
<< metal2 >>
rect -106 1542 1956 1598
rect -106 1478 -76 1542
rect 1916 1478 1956 1542
rect -106 1470 1956 1478
rect 30 1220 94 1226
rect 30 1214 36 1220
rect 88 1214 94 1220
rect 30 802 34 1214
rect 90 802 94 1214
rect 30 798 36 802
rect 88 798 94 802
rect 30 792 94 798
rect 124 1224 188 1470
rect 124 798 130 1224
rect 182 798 188 1224
rect 30 542 94 548
rect 30 536 36 542
rect 88 536 94 542
rect 30 124 34 536
rect 90 124 94 536
rect 30 120 36 124
rect 88 120 94 124
rect 30 114 94 120
rect 124 546 188 798
rect 222 1220 286 1226
rect 222 1214 228 1220
rect 280 1214 286 1220
rect 222 802 226 1214
rect 282 802 286 1214
rect 222 798 228 802
rect 280 798 286 802
rect 222 792 286 798
rect 316 1224 380 1470
rect 508 1462 1242 1470
rect 316 798 322 1224
rect 374 798 380 1224
rect 124 120 130 546
rect 182 120 188 546
rect 124 114 188 120
rect 222 542 286 548
rect 222 536 228 542
rect 280 536 286 542
rect 222 124 226 536
rect 282 124 286 536
rect 222 120 228 124
rect 280 120 286 124
rect 222 114 286 120
rect 316 546 380 798
rect 414 1220 478 1226
rect 414 1214 420 1220
rect 472 1214 478 1220
rect 414 802 418 1214
rect 474 802 478 1214
rect 414 798 420 802
rect 472 798 478 802
rect 414 792 478 798
rect 508 1224 572 1462
rect 508 798 514 1224
rect 566 798 572 1224
rect 316 120 322 546
rect 374 120 380 546
rect 316 114 380 120
rect 414 542 478 548
rect 414 536 420 542
rect 472 536 478 542
rect 414 124 418 536
rect 474 124 478 536
rect 414 120 420 124
rect 472 120 478 124
rect 414 114 478 120
rect 508 546 572 798
rect 606 1220 670 1226
rect 606 1214 612 1220
rect 664 1214 670 1220
rect 606 802 610 1214
rect 666 802 670 1214
rect 606 798 612 802
rect 664 798 670 802
rect 606 792 670 798
rect 700 1224 764 1462
rect 700 798 706 1224
rect 758 798 764 1224
rect 508 120 514 546
rect 566 120 572 546
rect 508 114 572 120
rect 606 542 670 548
rect 606 536 612 542
rect 664 536 670 542
rect 606 124 610 536
rect 666 124 670 536
rect 606 120 612 124
rect 664 120 670 124
rect 606 114 670 120
rect 700 546 764 798
rect 798 1220 862 1226
rect 798 1214 804 1220
rect 856 1214 862 1220
rect 798 802 802 1214
rect 858 802 862 1214
rect 798 798 804 802
rect 856 798 862 802
rect 798 792 862 798
rect 892 1224 956 1462
rect 892 798 898 1224
rect 950 798 956 1224
rect 700 120 706 546
rect 758 120 764 546
rect 700 114 764 120
rect 798 542 862 548
rect 798 536 804 542
rect 856 536 862 542
rect 798 124 802 536
rect 858 124 862 536
rect 798 120 804 124
rect 856 120 862 124
rect 798 114 862 120
rect 892 546 956 798
rect 990 1220 1054 1226
rect 990 1214 996 1220
rect 1048 1214 1054 1220
rect 990 802 994 1214
rect 1050 802 1054 1214
rect 990 798 996 802
rect 1048 798 1054 802
rect 990 792 1054 798
rect 1084 1224 1148 1462
rect 1084 798 1090 1224
rect 1142 798 1148 1224
rect 892 120 898 546
rect 950 120 956 546
rect 892 114 956 120
rect 990 542 1054 548
rect 990 536 996 542
rect 1048 536 1054 542
rect 990 124 994 536
rect 1050 124 1054 536
rect 990 120 996 124
rect 1048 120 1054 124
rect 990 114 1054 120
rect 1084 546 1148 798
rect 1182 1220 1246 1226
rect 1182 1214 1188 1220
rect 1240 1214 1246 1220
rect 1182 802 1186 1214
rect 1242 802 1246 1214
rect 1182 798 1188 802
rect 1240 798 1246 802
rect 1182 792 1246 798
rect 1276 1224 1340 1470
rect 1276 798 1282 1224
rect 1334 798 1340 1224
rect 1084 120 1090 546
rect 1142 120 1148 546
rect 1084 114 1148 120
rect 1182 542 1246 548
rect 1182 536 1188 542
rect 1240 536 1246 542
rect 1182 124 1186 536
rect 1242 124 1246 536
rect 1182 120 1188 124
rect 1240 120 1246 124
rect 1182 114 1246 120
rect 1276 546 1340 798
rect 1374 1220 1438 1226
rect 1374 1214 1380 1220
rect 1432 1214 1438 1220
rect 1374 802 1378 1214
rect 1434 802 1438 1214
rect 1374 798 1380 802
rect 1432 798 1438 802
rect 1374 792 1438 798
rect 1468 1224 1532 1470
rect 1468 798 1474 1224
rect 1526 798 1532 1224
rect 1276 120 1282 546
rect 1334 120 1340 546
rect 1276 114 1340 120
rect 1374 542 1438 548
rect 1374 536 1380 542
rect 1432 536 1438 542
rect 1374 124 1378 536
rect 1434 124 1438 536
rect 1374 120 1380 124
rect 1432 120 1438 124
rect 1374 114 1438 120
rect 1468 546 1532 798
rect 1566 1220 1630 1226
rect 1566 1214 1572 1220
rect 1624 1214 1630 1220
rect 1566 802 1570 1214
rect 1626 802 1630 1214
rect 1566 798 1572 802
rect 1624 798 1630 802
rect 1566 792 1630 798
rect 1660 1224 1724 1470
rect 1660 798 1666 1224
rect 1718 798 1724 1224
rect 1468 120 1474 546
rect 1526 120 1532 546
rect 1468 114 1532 120
rect 1566 542 1630 548
rect 1566 536 1572 542
rect 1624 536 1630 542
rect 1566 124 1570 536
rect 1626 124 1630 536
rect 1566 120 1572 124
rect 1624 120 1630 124
rect 1566 114 1630 120
rect 1660 546 1724 798
rect 1758 1220 1822 1226
rect 1758 1214 1764 1220
rect 1816 1214 1822 1220
rect 1758 802 1762 1214
rect 1818 802 1822 1214
rect 1758 798 1764 802
rect 1816 798 1822 802
rect 1758 792 1822 798
rect 1660 120 1666 546
rect 1718 120 1724 546
rect 1660 114 1724 120
rect 1758 542 1822 548
rect 1758 536 1764 542
rect 1816 536 1822 542
rect 1758 124 1762 536
rect 1818 124 1822 536
rect 1758 120 1764 124
rect 1816 120 1822 124
rect 1758 114 1822 120
rect 34 -350 100 -342
rect 34 -352 40 -350
rect 92 -352 100 -350
rect 34 -524 38 -352
rect 94 -524 100 -352
rect 34 -526 40 -524
rect 92 -526 100 -524
rect 34 -534 100 -526
rect 130 -350 194 -344
rect 130 -524 136 -350
rect 188 -524 194 -350
rect 34 -758 100 -750
rect 34 -760 40 -758
rect 92 -760 100 -758
rect 34 -932 38 -760
rect 94 -932 100 -760
rect 34 -934 40 -932
rect 92 -934 100 -932
rect 34 -942 100 -934
rect 130 -760 194 -524
rect 226 -350 292 -342
rect 226 -352 232 -350
rect 284 -352 292 -350
rect 226 -524 230 -352
rect 286 -524 292 -352
rect 226 -526 232 -524
rect 284 -526 292 -524
rect 226 -534 292 -526
rect 322 -350 386 -344
rect 322 -524 328 -350
rect 380 -524 386 -350
rect 130 -934 136 -760
rect 188 -934 194 -760
rect 130 -1142 194 -934
rect 226 -758 292 -750
rect 226 -760 232 -758
rect 284 -760 292 -758
rect 226 -932 230 -760
rect 286 -932 292 -760
rect 226 -934 232 -932
rect 284 -934 292 -932
rect 226 -942 292 -934
rect 322 -760 386 -524
rect 418 -350 484 -342
rect 418 -352 424 -350
rect 476 -352 484 -350
rect 418 -524 422 -352
rect 478 -524 484 -352
rect 418 -526 424 -524
rect 476 -526 484 -524
rect 418 -534 484 -526
rect 514 -350 578 -344
rect 514 -524 520 -350
rect 572 -524 578 -350
rect 322 -934 328 -760
rect 380 -934 386 -760
rect 322 -1142 386 -934
rect 418 -758 484 -750
rect 418 -760 424 -758
rect 476 -760 484 -758
rect 418 -932 422 -760
rect 478 -932 484 -760
rect 418 -934 424 -932
rect 476 -934 484 -932
rect 418 -942 484 -934
rect 514 -760 578 -524
rect 610 -350 676 -342
rect 610 -352 616 -350
rect 668 -352 676 -350
rect 610 -524 614 -352
rect 670 -524 676 -352
rect 610 -526 616 -524
rect 668 -526 676 -524
rect 610 -534 676 -526
rect 706 -350 770 -344
rect 706 -524 712 -350
rect 764 -524 770 -350
rect 514 -934 520 -760
rect 572 -934 578 -760
rect 514 -1142 578 -934
rect 610 -758 676 -750
rect 610 -760 616 -758
rect 668 -760 676 -758
rect 610 -932 614 -760
rect 670 -932 676 -760
rect 610 -934 616 -932
rect 668 -934 676 -932
rect 610 -942 676 -934
rect 706 -760 770 -524
rect 802 -350 868 -342
rect 802 -352 808 -350
rect 860 -352 868 -350
rect 802 -524 806 -352
rect 862 -524 868 -352
rect 802 -526 808 -524
rect 860 -526 868 -524
rect 802 -534 868 -526
rect 898 -350 962 -344
rect 898 -524 904 -350
rect 956 -524 962 -350
rect 706 -934 712 -760
rect 764 -934 770 -760
rect 706 -1142 770 -934
rect 802 -758 868 -750
rect 802 -760 808 -758
rect 860 -760 868 -758
rect 802 -932 806 -760
rect 862 -932 868 -760
rect 802 -934 808 -932
rect 860 -934 868 -932
rect 802 -942 868 -934
rect 898 -760 962 -524
rect 994 -350 1060 -342
rect 994 -352 1000 -350
rect 1052 -352 1060 -350
rect 994 -524 998 -352
rect 1054 -524 1060 -352
rect 994 -526 1000 -524
rect 1052 -526 1060 -524
rect 994 -534 1060 -526
rect 1090 -350 1154 -344
rect 1090 -524 1096 -350
rect 1148 -524 1154 -350
rect 898 -934 904 -760
rect 956 -934 962 -760
rect 898 -1142 962 -934
rect 994 -758 1060 -750
rect 994 -760 1000 -758
rect 1052 -760 1060 -758
rect 994 -932 998 -760
rect 1054 -932 1060 -760
rect 994 -934 1000 -932
rect 1052 -934 1060 -932
rect 994 -942 1060 -934
rect 1090 -760 1154 -524
rect 1186 -350 1252 -342
rect 1186 -352 1192 -350
rect 1244 -352 1252 -350
rect 1186 -524 1190 -352
rect 1246 -524 1252 -352
rect 1186 -526 1192 -524
rect 1244 -526 1252 -524
rect 1186 -534 1252 -526
rect 1282 -350 1346 -344
rect 1282 -524 1288 -350
rect 1340 -524 1346 -350
rect 1090 -934 1096 -760
rect 1148 -934 1154 -760
rect 1090 -1142 1154 -934
rect 1186 -758 1252 -750
rect 1186 -760 1192 -758
rect 1244 -760 1252 -758
rect 1186 -932 1190 -760
rect 1246 -932 1252 -760
rect 1186 -934 1192 -932
rect 1244 -934 1252 -932
rect 1186 -942 1252 -934
rect 1282 -760 1346 -524
rect 1378 -350 1444 -342
rect 1378 -352 1384 -350
rect 1436 -352 1444 -350
rect 1378 -524 1382 -352
rect 1438 -524 1444 -352
rect 1378 -526 1384 -524
rect 1436 -526 1444 -524
rect 1378 -534 1444 -526
rect 1474 -350 1538 -344
rect 1474 -524 1480 -350
rect 1532 -524 1538 -350
rect 1282 -934 1288 -760
rect 1340 -934 1346 -760
rect 1282 -1142 1346 -934
rect 1378 -758 1444 -750
rect 1378 -760 1384 -758
rect 1436 -760 1444 -758
rect 1378 -932 1382 -760
rect 1438 -932 1444 -760
rect 1378 -934 1384 -932
rect 1436 -934 1444 -932
rect 1378 -942 1444 -934
rect 1474 -760 1538 -524
rect 1570 -350 1636 -342
rect 1570 -352 1576 -350
rect 1628 -352 1636 -350
rect 1570 -524 1574 -352
rect 1630 -524 1636 -352
rect 1570 -526 1576 -524
rect 1628 -526 1636 -524
rect 1570 -534 1636 -526
rect 1666 -350 1730 -344
rect 1666 -524 1672 -350
rect 1724 -524 1730 -350
rect 1474 -934 1480 -760
rect 1532 -934 1538 -760
rect 1474 -1142 1538 -934
rect 1570 -758 1636 -750
rect 1570 -760 1576 -758
rect 1628 -760 1636 -758
rect 1570 -932 1574 -760
rect 1630 -932 1636 -760
rect 1570 -934 1576 -932
rect 1628 -934 1636 -932
rect 1570 -942 1636 -934
rect 1666 -760 1730 -524
rect 1762 -350 1828 -342
rect 1762 -352 1768 -350
rect 1820 -352 1828 -350
rect 1762 -524 1766 -352
rect 1822 -524 1828 -352
rect 1762 -526 1768 -524
rect 1820 -526 1828 -524
rect 1762 -534 1828 -526
rect 1666 -934 1672 -760
rect 1724 -934 1730 -760
rect 1666 -1142 1730 -934
rect 1762 -758 1828 -750
rect 1762 -760 1768 -758
rect 1820 -760 1828 -758
rect 1762 -932 1766 -760
rect 1822 -932 1828 -760
rect 1762 -934 1768 -932
rect 1820 -934 1828 -932
rect 1762 -942 1828 -934
rect -84 -1150 1940 -1142
rect -84 -1164 -64 -1150
rect -104 -1238 -64 -1164
rect 1922 -1164 1940 -1150
rect 1922 -1238 1958 -1164
rect -104 -1292 1958 -1238
<< via2 >>
rect 34 802 36 1214
rect 36 802 88 1214
rect 88 802 90 1214
rect 34 124 36 536
rect 36 124 88 536
rect 88 124 90 536
rect 226 802 228 1214
rect 228 802 280 1214
rect 280 802 282 1214
rect 226 124 228 536
rect 228 124 280 536
rect 280 124 282 536
rect 418 802 420 1214
rect 420 802 472 1214
rect 472 802 474 1214
rect 418 124 420 536
rect 420 124 472 536
rect 472 124 474 536
rect 610 802 612 1214
rect 612 802 664 1214
rect 664 802 666 1214
rect 610 124 612 536
rect 612 124 664 536
rect 664 124 666 536
rect 802 802 804 1214
rect 804 802 856 1214
rect 856 802 858 1214
rect 802 124 804 536
rect 804 124 856 536
rect 856 124 858 536
rect 994 802 996 1214
rect 996 802 1048 1214
rect 1048 802 1050 1214
rect 994 124 996 536
rect 996 124 1048 536
rect 1048 124 1050 536
rect 1186 802 1188 1214
rect 1188 802 1240 1214
rect 1240 802 1242 1214
rect 1186 124 1188 536
rect 1188 124 1240 536
rect 1240 124 1242 536
rect 1378 802 1380 1214
rect 1380 802 1432 1214
rect 1432 802 1434 1214
rect 1378 124 1380 536
rect 1380 124 1432 536
rect 1432 124 1434 536
rect 1570 802 1572 1214
rect 1572 802 1624 1214
rect 1624 802 1626 1214
rect 1570 124 1572 536
rect 1572 124 1624 536
rect 1624 124 1626 536
rect 1762 802 1764 1214
rect 1764 802 1816 1214
rect 1816 802 1818 1214
rect 1762 124 1764 536
rect 1764 124 1816 536
rect 1816 124 1818 536
rect 38 -524 40 -352
rect 40 -524 92 -352
rect 92 -524 94 -352
rect 38 -932 40 -760
rect 40 -932 92 -760
rect 92 -932 94 -760
rect 230 -524 232 -352
rect 232 -524 284 -352
rect 284 -524 286 -352
rect 230 -932 232 -760
rect 232 -932 284 -760
rect 284 -932 286 -760
rect 422 -524 424 -352
rect 424 -524 476 -352
rect 476 -524 478 -352
rect 422 -932 424 -760
rect 424 -932 476 -760
rect 476 -932 478 -760
rect 614 -524 616 -352
rect 616 -524 668 -352
rect 668 -524 670 -352
rect 614 -932 616 -760
rect 616 -932 668 -760
rect 668 -932 670 -760
rect 806 -524 808 -352
rect 808 -524 860 -352
rect 860 -524 862 -352
rect 806 -932 808 -760
rect 808 -932 860 -760
rect 860 -932 862 -760
rect 998 -524 1000 -352
rect 1000 -524 1052 -352
rect 1052 -524 1054 -352
rect 998 -932 1000 -760
rect 1000 -932 1052 -760
rect 1052 -932 1054 -760
rect 1190 -524 1192 -352
rect 1192 -524 1244 -352
rect 1244 -524 1246 -352
rect 1190 -932 1192 -760
rect 1192 -932 1244 -760
rect 1244 -932 1246 -760
rect 1382 -524 1384 -352
rect 1384 -524 1436 -352
rect 1436 -524 1438 -352
rect 1382 -932 1384 -760
rect 1384 -932 1436 -760
rect 1436 -932 1438 -760
rect 1574 -524 1576 -352
rect 1576 -524 1628 -352
rect 1628 -524 1630 -352
rect 1574 -932 1576 -760
rect 1576 -932 1628 -760
rect 1628 -932 1630 -760
rect 1766 -524 1768 -352
rect 1768 -524 1820 -352
rect 1820 -524 1822 -352
rect 1766 -932 1768 -760
rect 1768 -932 1820 -760
rect 1820 -932 1822 -760
<< metal3 >>
rect 28 1214 96 1228
rect 28 802 34 1214
rect 90 802 96 1214
rect 28 536 96 802
rect 28 124 34 536
rect 90 124 96 536
rect 28 -36 96 124
rect 220 1214 288 1228
rect 220 802 226 1214
rect 282 802 288 1214
rect 220 536 288 802
rect 220 124 226 536
rect 282 124 288 536
rect 220 -36 288 124
rect 412 1214 480 1228
rect 412 802 418 1214
rect 474 802 480 1214
rect 412 536 480 802
rect 412 124 418 536
rect 474 124 480 536
rect 412 -36 480 124
rect 604 1214 672 1228
rect 604 802 610 1214
rect 666 802 672 1214
rect 604 536 672 802
rect 604 124 610 536
rect 666 124 672 536
rect 604 -36 672 124
rect 796 1214 864 1228
rect 796 802 802 1214
rect 858 802 864 1214
rect 796 536 864 802
rect 796 124 802 536
rect 858 124 864 536
rect 796 -36 864 124
rect 988 1214 1056 1228
rect 988 802 994 1214
rect 1050 802 1056 1214
rect 988 536 1056 802
rect 988 124 994 536
rect 1050 124 1056 536
rect 988 -36 1056 124
rect 1180 1214 1248 1228
rect 1180 802 1186 1214
rect 1242 802 1248 1214
rect 1180 536 1248 802
rect 1180 124 1186 536
rect 1242 124 1248 536
rect 1180 -36 1248 124
rect 1372 1214 1440 1228
rect 1372 802 1378 1214
rect 1434 802 1440 1214
rect 1372 536 1440 802
rect 1372 124 1378 536
rect 1434 124 1440 536
rect 1372 -36 1440 124
rect 1564 1214 1632 1228
rect 1564 802 1570 1214
rect 1626 802 1632 1214
rect 1564 536 1632 802
rect 1564 124 1570 536
rect 1626 124 1632 536
rect 1564 -36 1632 124
rect 1756 1214 1824 1228
rect 1756 802 1762 1214
rect 1818 802 1824 1214
rect 1756 536 1824 802
rect 1756 124 1762 536
rect 1818 124 1824 536
rect 1756 -36 1824 124
rect 28 -200 1986 -36
rect 32 -352 100 -200
rect 32 -524 38 -352
rect 94 -524 100 -352
rect 32 -760 100 -524
rect 32 -932 38 -760
rect 94 -932 100 -760
rect 32 -942 100 -932
rect 224 -352 292 -200
rect 224 -524 230 -352
rect 286 -524 292 -352
rect 224 -760 292 -524
rect 224 -932 230 -760
rect 286 -932 292 -760
rect 224 -942 292 -932
rect 416 -352 484 -200
rect 416 -524 422 -352
rect 478 -524 484 -352
rect 416 -760 484 -524
rect 416 -932 422 -760
rect 478 -932 484 -760
rect 416 -942 484 -932
rect 608 -352 676 -200
rect 608 -524 614 -352
rect 670 -524 676 -352
rect 608 -760 676 -524
rect 608 -932 614 -760
rect 670 -932 676 -760
rect 608 -942 676 -932
rect 800 -352 868 -200
rect 800 -524 806 -352
rect 862 -524 868 -352
rect 800 -760 868 -524
rect 800 -932 806 -760
rect 862 -932 868 -760
rect 800 -942 868 -932
rect 992 -352 1060 -200
rect 992 -524 998 -352
rect 1054 -524 1060 -352
rect 992 -760 1060 -524
rect 992 -932 998 -760
rect 1054 -932 1060 -760
rect 992 -942 1060 -932
rect 1184 -352 1252 -200
rect 1184 -524 1190 -352
rect 1246 -524 1252 -352
rect 1184 -760 1252 -524
rect 1184 -932 1190 -760
rect 1246 -932 1252 -760
rect 1184 -942 1252 -932
rect 1376 -352 1444 -200
rect 1376 -524 1382 -352
rect 1438 -524 1444 -352
rect 1376 -760 1444 -524
rect 1376 -932 1382 -760
rect 1438 -932 1444 -760
rect 1376 -942 1444 -932
rect 1568 -352 1636 -200
rect 1568 -524 1574 -352
rect 1630 -524 1636 -352
rect 1568 -760 1636 -524
rect 1568 -932 1574 -760
rect 1630 -932 1636 -760
rect 1568 -942 1636 -932
rect 1760 -352 1828 -200
rect 1760 -524 1766 -352
rect 1822 -524 1828 -352
rect 1760 -760 1828 -524
rect 1760 -932 1766 -760
rect 1822 -932 1828 -760
rect 1760 -942 1828 -932
use sky130_fd_pr__pfet_01v8_VNEHM9  sky130_fd_pr__pfet_01v8_VNEHM9_0
timestamp 1627668659
transform 1 0 925 0 1 673
box -1031 -779 1031 779
use sky130_fd_pr__nfet_01v8_BBTBMZ  sky130_fd_pr__nfet_01v8_BBTBMZ_0
timestamp 1627668659
transform 1 0 929 0 1 -641
box -1031 -511 1031 511
<< labels >>
rlabel metal3 1934 -200 1986 -36 1 out
port 3 n
rlabel metal2 -100 1480 1946 1582 1 VDD
port 4 n
rlabel metal2 -94 -1278 1952 -1176 1 GND
port 2 n
rlabel metal1 -160 -220 -16 -16 1 in
port 5 n
<< end >>
