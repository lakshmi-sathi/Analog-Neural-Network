magic
tech sky130A
magscale 1 2
timestamp 1628060682
<< error_p >>
rect -749 549 -691 555
rect -557 549 -499 555
rect -365 549 -307 555
rect -173 549 -115 555
rect 19 549 77 555
rect 211 549 269 555
rect 403 549 461 555
rect 595 549 653 555
rect -749 515 -737 549
rect -557 515 -545 549
rect -365 515 -353 549
rect -173 515 -161 549
rect 19 515 31 549
rect 211 515 223 549
rect 403 515 415 549
rect 595 515 607 549
rect -749 509 -691 515
rect -557 509 -499 515
rect -365 509 -307 515
rect -173 509 -115 515
rect 19 509 77 515
rect 211 509 269 515
rect 403 509 461 515
rect 595 509 653 515
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect -749 -515 -691 -509
rect -557 -515 -499 -509
rect -365 -515 -307 -509
rect -173 -515 -115 -509
rect 19 -515 77 -509
rect 211 -515 269 -509
rect 403 -515 461 -509
rect 595 -515 653 -509
rect -749 -549 -737 -515
rect -557 -549 -545 -515
rect -365 -549 -353 -515
rect -173 -549 -161 -515
rect 19 -549 31 -515
rect 211 -549 223 -515
rect 403 -549 415 -515
rect 595 -549 607 -515
rect -749 -555 -691 -549
rect -557 -555 -499 -549
rect -365 -555 -307 -549
rect -173 -555 -115 -549
rect 19 -555 77 -549
rect 211 -555 269 -549
rect 403 -555 461 -549
rect 595 -555 653 -549
<< nwell >>
rect -935 -687 935 687
<< pmos >>
rect -735 118 -705 468
rect -639 118 -609 468
rect -543 118 -513 468
rect -447 118 -417 468
rect -351 118 -321 468
rect -255 118 -225 468
rect -159 118 -129 468
rect -63 118 -33 468
rect 33 118 63 468
rect 129 118 159 468
rect 225 118 255 468
rect 321 118 351 468
rect 417 118 447 468
rect 513 118 543 468
rect 609 118 639 468
rect 705 118 735 468
rect -735 -468 -705 -118
rect -639 -468 -609 -118
rect -543 -468 -513 -118
rect -447 -468 -417 -118
rect -351 -468 -321 -118
rect -255 -468 -225 -118
rect -159 -468 -129 -118
rect -63 -468 -33 -118
rect 33 -468 63 -118
rect 129 -468 159 -118
rect 225 -468 255 -118
rect 321 -468 351 -118
rect 417 -468 447 -118
rect 513 -468 543 -118
rect 609 -468 639 -118
rect 705 -468 735 -118
<< pdiff >>
rect -797 456 -735 468
rect -797 130 -785 456
rect -751 130 -735 456
rect -797 118 -735 130
rect -705 456 -639 468
rect -705 130 -689 456
rect -655 130 -639 456
rect -705 118 -639 130
rect -609 456 -543 468
rect -609 130 -593 456
rect -559 130 -543 456
rect -609 118 -543 130
rect -513 456 -447 468
rect -513 130 -497 456
rect -463 130 -447 456
rect -513 118 -447 130
rect -417 456 -351 468
rect -417 130 -401 456
rect -367 130 -351 456
rect -417 118 -351 130
rect -321 456 -255 468
rect -321 130 -305 456
rect -271 130 -255 456
rect -321 118 -255 130
rect -225 456 -159 468
rect -225 130 -209 456
rect -175 130 -159 456
rect -225 118 -159 130
rect -129 456 -63 468
rect -129 130 -113 456
rect -79 130 -63 456
rect -129 118 -63 130
rect -33 456 33 468
rect -33 130 -17 456
rect 17 130 33 456
rect -33 118 33 130
rect 63 456 129 468
rect 63 130 79 456
rect 113 130 129 456
rect 63 118 129 130
rect 159 456 225 468
rect 159 130 175 456
rect 209 130 225 456
rect 159 118 225 130
rect 255 456 321 468
rect 255 130 271 456
rect 305 130 321 456
rect 255 118 321 130
rect 351 456 417 468
rect 351 130 367 456
rect 401 130 417 456
rect 351 118 417 130
rect 447 456 513 468
rect 447 130 463 456
rect 497 130 513 456
rect 447 118 513 130
rect 543 456 609 468
rect 543 130 559 456
rect 593 130 609 456
rect 543 118 609 130
rect 639 456 705 468
rect 639 130 655 456
rect 689 130 705 456
rect 639 118 705 130
rect 735 456 797 468
rect 735 130 751 456
rect 785 130 797 456
rect 735 118 797 130
rect -797 -130 -735 -118
rect -797 -456 -785 -130
rect -751 -456 -735 -130
rect -797 -468 -735 -456
rect -705 -130 -639 -118
rect -705 -456 -689 -130
rect -655 -456 -639 -130
rect -705 -468 -639 -456
rect -609 -130 -543 -118
rect -609 -456 -593 -130
rect -559 -456 -543 -130
rect -609 -468 -543 -456
rect -513 -130 -447 -118
rect -513 -456 -497 -130
rect -463 -456 -447 -130
rect -513 -468 -447 -456
rect -417 -130 -351 -118
rect -417 -456 -401 -130
rect -367 -456 -351 -130
rect -417 -468 -351 -456
rect -321 -130 -255 -118
rect -321 -456 -305 -130
rect -271 -456 -255 -130
rect -321 -468 -255 -456
rect -225 -130 -159 -118
rect -225 -456 -209 -130
rect -175 -456 -159 -130
rect -225 -468 -159 -456
rect -129 -130 -63 -118
rect -129 -456 -113 -130
rect -79 -456 -63 -130
rect -129 -468 -63 -456
rect -33 -130 33 -118
rect -33 -456 -17 -130
rect 17 -456 33 -130
rect -33 -468 33 -456
rect 63 -130 129 -118
rect 63 -456 79 -130
rect 113 -456 129 -130
rect 63 -468 129 -456
rect 159 -130 225 -118
rect 159 -456 175 -130
rect 209 -456 225 -130
rect 159 -468 225 -456
rect 255 -130 321 -118
rect 255 -456 271 -130
rect 305 -456 321 -130
rect 255 -468 321 -456
rect 351 -130 417 -118
rect 351 -456 367 -130
rect 401 -456 417 -130
rect 351 -468 417 -456
rect 447 -130 513 -118
rect 447 -456 463 -130
rect 497 -456 513 -130
rect 447 -468 513 -456
rect 543 -130 609 -118
rect 543 -456 559 -130
rect 593 -456 609 -130
rect 543 -468 609 -456
rect 639 -130 705 -118
rect 639 -456 655 -130
rect 689 -456 705 -130
rect 639 -468 705 -456
rect 735 -130 797 -118
rect 735 -456 751 -130
rect 785 -456 797 -130
rect 735 -468 797 -456
<< pdiffc >>
rect -785 130 -751 456
rect -689 130 -655 456
rect -593 130 -559 456
rect -497 130 -463 456
rect -401 130 -367 456
rect -305 130 -271 456
rect -209 130 -175 456
rect -113 130 -79 456
rect -17 130 17 456
rect 79 130 113 456
rect 175 130 209 456
rect 271 130 305 456
rect 367 130 401 456
rect 463 130 497 456
rect 559 130 593 456
rect 655 130 689 456
rect 751 130 785 456
rect -785 -456 -751 -130
rect -689 -456 -655 -130
rect -593 -456 -559 -130
rect -497 -456 -463 -130
rect -401 -456 -367 -130
rect -305 -456 -271 -130
rect -209 -456 -175 -130
rect -113 -456 -79 -130
rect -17 -456 17 -130
rect 79 -456 113 -130
rect 175 -456 209 -130
rect 271 -456 305 -130
rect 367 -456 401 -130
rect 463 -456 497 -130
rect 559 -456 593 -130
rect 655 -456 689 -130
rect 751 -456 785 -130
<< nsubdiff >>
rect -899 617 -803 651
rect 803 617 899 651
rect -899 555 -865 617
rect 865 555 899 617
rect -899 -617 -865 -555
rect 865 -617 899 -555
rect -899 -651 -803 -617
rect 803 -651 899 -617
<< nsubdiffcont >>
rect -803 617 803 651
rect -899 -555 -865 555
rect 865 -555 899 555
rect -803 -651 803 -617
<< poly >>
rect -753 549 -687 565
rect -753 515 -737 549
rect -703 515 -687 549
rect -753 499 -687 515
rect -561 549 -495 565
rect -561 515 -545 549
rect -511 515 -495 549
rect -561 499 -495 515
rect -369 549 -303 565
rect -369 515 -353 549
rect -319 515 -303 549
rect -369 499 -303 515
rect -177 549 -111 565
rect -177 515 -161 549
rect -127 515 -111 549
rect -177 499 -111 515
rect 15 549 81 565
rect 15 515 31 549
rect 65 515 81 549
rect 15 499 81 515
rect 207 549 273 565
rect 207 515 223 549
rect 257 515 273 549
rect 207 499 273 515
rect 399 549 465 565
rect 399 515 415 549
rect 449 515 465 549
rect 399 499 465 515
rect 591 549 657 565
rect 591 515 607 549
rect 641 515 657 549
rect 591 499 657 515
rect -735 468 -705 499
rect -639 468 -609 494
rect -543 468 -513 499
rect -447 468 -417 494
rect -351 468 -321 499
rect -255 468 -225 494
rect -159 468 -129 499
rect -63 468 -33 494
rect 33 468 63 499
rect 129 468 159 494
rect 225 468 255 499
rect 321 468 351 494
rect 417 468 447 499
rect 513 468 543 494
rect 609 468 639 499
rect 705 468 735 494
rect -735 92 -705 118
rect -639 87 -609 118
rect -543 92 -513 118
rect -447 87 -417 118
rect -351 92 -321 118
rect -255 87 -225 118
rect -159 92 -129 118
rect -63 87 -33 118
rect 33 92 63 118
rect 129 87 159 118
rect 225 92 255 118
rect 321 87 351 118
rect 417 92 447 118
rect 513 87 543 118
rect 609 92 639 118
rect 705 87 735 118
rect -657 71 -591 87
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 687 -87 753 -71
rect -735 -118 -705 -92
rect -639 -118 -609 -87
rect -543 -118 -513 -92
rect -447 -118 -417 -87
rect -351 -118 -321 -92
rect -255 -118 -225 -87
rect -159 -118 -129 -92
rect -63 -118 -33 -87
rect 33 -118 63 -92
rect 129 -118 159 -87
rect 225 -118 255 -92
rect 321 -118 351 -87
rect 417 -118 447 -92
rect 513 -118 543 -87
rect 609 -118 639 -92
rect 705 -118 735 -87
rect -735 -499 -705 -468
rect -639 -494 -609 -468
rect -543 -499 -513 -468
rect -447 -494 -417 -468
rect -351 -499 -321 -468
rect -255 -494 -225 -468
rect -159 -499 -129 -468
rect -63 -494 -33 -468
rect 33 -499 63 -468
rect 129 -494 159 -468
rect 225 -499 255 -468
rect 321 -494 351 -468
rect 417 -499 447 -468
rect 513 -494 543 -468
rect 609 -499 639 -468
rect 705 -494 735 -468
rect -753 -515 -687 -499
rect -753 -549 -737 -515
rect -703 -549 -687 -515
rect -753 -565 -687 -549
rect -561 -515 -495 -499
rect -561 -549 -545 -515
rect -511 -549 -495 -515
rect -561 -565 -495 -549
rect -369 -515 -303 -499
rect -369 -549 -353 -515
rect -319 -549 -303 -515
rect -369 -565 -303 -549
rect -177 -515 -111 -499
rect -177 -549 -161 -515
rect -127 -549 -111 -515
rect -177 -565 -111 -549
rect 15 -515 81 -499
rect 15 -549 31 -515
rect 65 -549 81 -515
rect 15 -565 81 -549
rect 207 -515 273 -499
rect 207 -549 223 -515
rect 257 -549 273 -515
rect 207 -565 273 -549
rect 399 -515 465 -499
rect 399 -549 415 -515
rect 449 -549 465 -515
rect 399 -565 465 -549
rect 591 -515 657 -499
rect 591 -549 607 -515
rect 641 -549 657 -515
rect 591 -565 657 -549
<< polycont >>
rect -737 515 -703 549
rect -545 515 -511 549
rect -353 515 -319 549
rect -161 515 -127 549
rect 31 515 65 549
rect 223 515 257 549
rect 415 515 449 549
rect 607 515 641 549
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect -737 -549 -703 -515
rect -545 -549 -511 -515
rect -353 -549 -319 -515
rect -161 -549 -127 -515
rect 31 -549 65 -515
rect 223 -549 257 -515
rect 415 -549 449 -515
rect 607 -549 641 -515
<< locali >>
rect -899 617 -803 651
rect 803 617 899 651
rect -899 555 -865 617
rect 865 555 899 617
rect -753 515 -737 549
rect -703 515 -687 549
rect -561 515 -545 549
rect -511 515 -495 549
rect -369 515 -353 549
rect -319 515 -303 549
rect -177 515 -161 549
rect -127 515 -111 549
rect 15 515 31 549
rect 65 515 81 549
rect 207 515 223 549
rect 257 515 273 549
rect 399 515 415 549
rect 449 515 465 549
rect 591 515 607 549
rect 641 515 657 549
rect -785 456 -751 472
rect -785 114 -751 130
rect -689 456 -655 472
rect -689 114 -655 130
rect -593 456 -559 472
rect -593 114 -559 130
rect -497 456 -463 472
rect -497 114 -463 130
rect -401 456 -367 472
rect -401 114 -367 130
rect -305 456 -271 472
rect -305 114 -271 130
rect -209 456 -175 472
rect -209 114 -175 130
rect -113 456 -79 472
rect -113 114 -79 130
rect -17 456 17 472
rect -17 114 17 130
rect 79 456 113 472
rect 79 114 113 130
rect 175 456 209 472
rect 175 114 209 130
rect 271 456 305 472
rect 271 114 305 130
rect 367 456 401 472
rect 367 114 401 130
rect 463 456 497 472
rect 463 114 497 130
rect 559 456 593 472
rect 559 114 593 130
rect 655 456 689 472
rect 655 114 689 130
rect 751 456 785 472
rect 751 114 785 130
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect -785 -130 -751 -114
rect -785 -472 -751 -456
rect -689 -130 -655 -114
rect -689 -472 -655 -456
rect -593 -130 -559 -114
rect -593 -472 -559 -456
rect -497 -130 -463 -114
rect -497 -472 -463 -456
rect -401 -130 -367 -114
rect -401 -472 -367 -456
rect -305 -130 -271 -114
rect -305 -472 -271 -456
rect -209 -130 -175 -114
rect -209 -472 -175 -456
rect -113 -130 -79 -114
rect -113 -472 -79 -456
rect -17 -130 17 -114
rect -17 -472 17 -456
rect 79 -130 113 -114
rect 79 -472 113 -456
rect 175 -130 209 -114
rect 175 -472 209 -456
rect 271 -130 305 -114
rect 271 -472 305 -456
rect 367 -130 401 -114
rect 367 -472 401 -456
rect 463 -130 497 -114
rect 463 -472 497 -456
rect 559 -130 593 -114
rect 559 -472 593 -456
rect 655 -130 689 -114
rect 655 -472 689 -456
rect 751 -130 785 -114
rect 751 -472 785 -456
rect -753 -549 -737 -515
rect -703 -549 -687 -515
rect -561 -549 -545 -515
rect -511 -549 -495 -515
rect -369 -549 -353 -515
rect -319 -549 -303 -515
rect -177 -549 -161 -515
rect -127 -549 -111 -515
rect 15 -549 31 -515
rect 65 -549 81 -515
rect 207 -549 223 -515
rect 257 -549 273 -515
rect 399 -549 415 -515
rect 449 -549 465 -515
rect 591 -549 607 -515
rect 641 -549 657 -515
rect -899 -617 -865 -555
rect 865 -617 899 -555
rect -899 -651 -803 -617
rect 803 -651 899 -617
<< viali >>
rect -737 515 -703 549
rect -545 515 -511 549
rect -353 515 -319 549
rect -161 515 -127 549
rect 31 515 65 549
rect 223 515 257 549
rect 415 515 449 549
rect 607 515 641 549
rect -785 130 -751 456
rect -689 130 -655 456
rect -593 130 -559 456
rect -497 130 -463 456
rect -401 130 -367 456
rect -305 130 -271 456
rect -209 130 -175 456
rect -113 130 -79 456
rect -17 130 17 456
rect 79 130 113 456
rect 175 130 209 456
rect 271 130 305 456
rect 367 130 401 456
rect 463 130 497 456
rect 559 130 593 456
rect 655 130 689 456
rect 751 130 785 456
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect -785 -456 -751 -130
rect -689 -456 -655 -130
rect -593 -456 -559 -130
rect -497 -456 -463 -130
rect -401 -456 -367 -130
rect -305 -456 -271 -130
rect -209 -456 -175 -130
rect -113 -456 -79 -130
rect -17 -456 17 -130
rect 79 -456 113 -130
rect 175 -456 209 -130
rect 271 -456 305 -130
rect 367 -456 401 -130
rect 463 -456 497 -130
rect 559 -456 593 -130
rect 655 -456 689 -130
rect 751 -456 785 -130
rect -737 -549 -703 -515
rect -545 -549 -511 -515
rect -353 -549 -319 -515
rect -161 -549 -127 -515
rect 31 -549 65 -515
rect 223 -549 257 -515
rect 415 -549 449 -515
rect 607 -549 641 -515
<< metal1 >>
rect -749 549 -691 555
rect -749 515 -737 549
rect -703 515 -691 549
rect -749 509 -691 515
rect -557 549 -499 555
rect -557 515 -545 549
rect -511 515 -499 549
rect -557 509 -499 515
rect -365 549 -307 555
rect -365 515 -353 549
rect -319 515 -307 549
rect -365 509 -307 515
rect -173 549 -115 555
rect -173 515 -161 549
rect -127 515 -115 549
rect -173 509 -115 515
rect 19 549 77 555
rect 19 515 31 549
rect 65 515 77 549
rect 19 509 77 515
rect 211 549 269 555
rect 211 515 223 549
rect 257 515 269 549
rect 211 509 269 515
rect 403 549 461 555
rect 403 515 415 549
rect 449 515 461 549
rect 403 509 461 515
rect 595 549 653 555
rect 595 515 607 549
rect 641 515 653 549
rect 595 509 653 515
rect -791 456 -745 468
rect -791 130 -785 456
rect -751 130 -745 456
rect -791 118 -745 130
rect -695 456 -649 468
rect -695 130 -689 456
rect -655 130 -649 456
rect -695 118 -649 130
rect -599 456 -553 468
rect -599 130 -593 456
rect -559 130 -553 456
rect -599 118 -553 130
rect -503 456 -457 468
rect -503 130 -497 456
rect -463 130 -457 456
rect -503 118 -457 130
rect -407 456 -361 468
rect -407 130 -401 456
rect -367 130 -361 456
rect -407 118 -361 130
rect -311 456 -265 468
rect -311 130 -305 456
rect -271 130 -265 456
rect -311 118 -265 130
rect -215 456 -169 468
rect -215 130 -209 456
rect -175 130 -169 456
rect -215 118 -169 130
rect -119 456 -73 468
rect -119 130 -113 456
rect -79 130 -73 456
rect -119 118 -73 130
rect -23 456 23 468
rect -23 130 -17 456
rect 17 130 23 456
rect -23 118 23 130
rect 73 456 119 468
rect 73 130 79 456
rect 113 130 119 456
rect 73 118 119 130
rect 169 456 215 468
rect 169 130 175 456
rect 209 130 215 456
rect 169 118 215 130
rect 265 456 311 468
rect 265 130 271 456
rect 305 130 311 456
rect 265 118 311 130
rect 361 456 407 468
rect 361 130 367 456
rect 401 130 407 456
rect 361 118 407 130
rect 457 456 503 468
rect 457 130 463 456
rect 497 130 503 456
rect 457 118 503 130
rect 553 456 599 468
rect 553 130 559 456
rect 593 130 599 456
rect 553 118 599 130
rect 649 456 695 468
rect 649 130 655 456
rect 689 130 695 456
rect 649 118 695 130
rect 745 456 791 468
rect 745 130 751 456
rect 785 130 791 456
rect 745 118 791 130
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect -791 -130 -745 -118
rect -791 -456 -785 -130
rect -751 -456 -745 -130
rect -791 -468 -745 -456
rect -695 -130 -649 -118
rect -695 -456 -689 -130
rect -655 -456 -649 -130
rect -695 -468 -649 -456
rect -599 -130 -553 -118
rect -599 -456 -593 -130
rect -559 -456 -553 -130
rect -599 -468 -553 -456
rect -503 -130 -457 -118
rect -503 -456 -497 -130
rect -463 -456 -457 -130
rect -503 -468 -457 -456
rect -407 -130 -361 -118
rect -407 -456 -401 -130
rect -367 -456 -361 -130
rect -407 -468 -361 -456
rect -311 -130 -265 -118
rect -311 -456 -305 -130
rect -271 -456 -265 -130
rect -311 -468 -265 -456
rect -215 -130 -169 -118
rect -215 -456 -209 -130
rect -175 -456 -169 -130
rect -215 -468 -169 -456
rect -119 -130 -73 -118
rect -119 -456 -113 -130
rect -79 -456 -73 -130
rect -119 -468 -73 -456
rect -23 -130 23 -118
rect -23 -456 -17 -130
rect 17 -456 23 -130
rect -23 -468 23 -456
rect 73 -130 119 -118
rect 73 -456 79 -130
rect 113 -456 119 -130
rect 73 -468 119 -456
rect 169 -130 215 -118
rect 169 -456 175 -130
rect 209 -456 215 -130
rect 169 -468 215 -456
rect 265 -130 311 -118
rect 265 -456 271 -130
rect 305 -456 311 -130
rect 265 -468 311 -456
rect 361 -130 407 -118
rect 361 -456 367 -130
rect 401 -456 407 -130
rect 361 -468 407 -456
rect 457 -130 503 -118
rect 457 -456 463 -130
rect 497 -456 503 -130
rect 457 -468 503 -456
rect 553 -130 599 -118
rect 553 -456 559 -130
rect 593 -456 599 -130
rect 553 -468 599 -456
rect 649 -130 695 -118
rect 649 -456 655 -130
rect 689 -456 695 -130
rect 649 -468 695 -456
rect 745 -130 791 -118
rect 745 -456 751 -130
rect 785 -456 791 -130
rect 745 -468 791 -456
rect -749 -515 -691 -509
rect -749 -549 -737 -515
rect -703 -549 -691 -515
rect -749 -555 -691 -549
rect -557 -515 -499 -509
rect -557 -549 -545 -515
rect -511 -549 -499 -515
rect -557 -555 -499 -549
rect -365 -515 -307 -509
rect -365 -549 -353 -515
rect -319 -549 -307 -515
rect -365 -555 -307 -549
rect -173 -515 -115 -509
rect -173 -549 -161 -515
rect -127 -549 -115 -515
rect -173 -555 -115 -549
rect 19 -515 77 -509
rect 19 -549 31 -515
rect 65 -549 77 -515
rect 19 -555 77 -549
rect 211 -515 269 -509
rect 211 -549 223 -515
rect 257 -549 269 -515
rect 211 -555 269 -549
rect 403 -515 461 -509
rect 403 -549 415 -515
rect 449 -549 461 -515
rect 403 -555 461 -549
rect 595 -515 653 -509
rect 595 -549 607 -515
rect 641 -549 653 -515
rect 595 -555 653 -549
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -882 -634 882 634
string parameters w 1.75 l 0.15 m 2 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
