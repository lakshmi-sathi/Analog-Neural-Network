magic
tech sky130A
magscale 1 2
timestamp 1628069922
<< xpolycontact >>
rect -69 95 69 527
rect -69 -527 69 -95
<< ppolyres >>
rect -69 -95 69 95
<< viali >>
rect -53 112 53 509
rect -53 -509 53 -112
<< metal1 >>
rect -59 509 59 521
rect -59 112 -53 509
rect 53 112 59 509
rect -59 100 59 112
rect -59 -112 59 -100
rect -59 -509 -53 -112
rect 53 -509 59 -112
rect -59 -521 59 -509
<< res0p69 >>
rect -71 -97 71 97
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p69
string parameters w 0.690 l 0.95 m 1 nx 1 wmin 0.690 lmin 0.50 rho 319.8 val 495.921 dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 0.690 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
