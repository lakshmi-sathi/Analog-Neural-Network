magic
tech sky130A
magscale 1 2
timestamp 1628105024
<< metal1 >>
rect -6183 4348 -4726 4674
rect -6176 1604 -4518 1896
rect 442 1736 1162 1752
rect 436 1270 446 1736
rect 1142 1270 1162 1736
rect 442 1210 1162 1270
rect 11910 1040 12486 1410
rect -6200 -1284 -4518 -992
<< via1 >>
rect 446 1270 1142 1736
<< metal2 >>
rect -2211 5291 -2105 5305
rect -2985 5275 -2387 5277
rect -2309 5275 -2105 5291
rect -2985 5171 -2105 5275
rect -2471 3445 -2105 5171
rect -2471 3326 12017 3445
rect -5430 2950 -4336 3074
rect -2471 3014 12020 3326
rect -5430 302 -5022 2950
rect -2471 2505 -2105 3014
rect -2929 2399 -2105 2505
rect -5430 178 -4424 302
rect -5430 -2578 -5022 178
rect -2471 -375 -2105 2399
rect 446 1736 1142 1746
rect 446 1260 1142 1270
rect 2042 98 2248 130
rect 1648 -290 11828 98
rect -2973 -481 -2105 -375
rect 2042 -2578 2430 -290
rect -5430 -2634 -4358 -2578
rect -3050 -2634 2430 -2578
rect -5494 -3042 2432 -2634
<< via2 >>
rect 446 1270 1142 1736
<< metal3 >>
rect -2651 3897 -2380 5933
rect -3113 3807 -2380 3897
rect -2033 1125 -1673 5938
rect -3049 1035 -1673 1125
rect -1209 -1755 -711 5957
rect 446 1741 1072 5990
rect 436 1736 1152 1741
rect 436 1270 446 1736
rect 1142 1270 1152 1736
rect 436 1265 1152 1270
rect 11886 190 13048 498
rect -3039 -1845 -711 -1755
use analogneuron_invopamp_re_15kfeedbck  analogneuron_invopamp_re_15kfeedbck_0
timestamp 1628105024
transform 1 0 1354 0 1 234
box -1354 -234 10724 2910
use aninv_  aninv__0
timestamp 1628080314
transform -1 0 -2858 0 1 3671
box -63 -721 1952 1584
use aninv_  aninv__1
timestamp 1628080314
transform -1 0 -2858 0 1 899
box -63 -721 1952 1584
use aninv_  aninv__2
timestamp 1628080314
transform -1 0 -2858 0 1 -1981
box -63 -721 1952 1584
<< labels >>
rlabel metal3 12386 200 13016 482 1 Out
port 1 n
rlabel metal1 -6158 4352 -5796 4664 1 In1
port 3 n
rlabel metal1 12116 1056 12472 1404 1 Vref
port 4 n
rlabel metal1 -6164 1612 -5830 1880 1 In2
port 5 n
rlabel metal1 -6176 -1274 -5842 -1006 1 In3
port 6 n
rlabel metal3 -2636 5770 -2388 5924 1 R1
port 7 n
rlabel metal3 -2018 5770 -1686 5926 1 R2
port 8 n
rlabel metal3 -1192 5782 -728 5942 1 R3
port 9 n
rlabel metal3 470 5766 1042 5966 1 amp_in
port 10 n
rlabel metal2 1706 3070 11834 3360 1 VDD
port 11 n
rlabel metal2 1726 -248 11738 2 1 GND
port 12 n
<< end >>
