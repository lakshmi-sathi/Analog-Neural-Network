magic
tech sky130A
magscale 1 2
timestamp 1627922418
<< xpolycontact >>
rect -35 295 35 727
rect -35 -727 35 -295
<< ppolyres >>
rect -35 -295 35 295
<< viali >>
rect -19 312 19 709
rect -19 -709 19 -312
<< metal1 >>
rect -25 709 25 721
rect -25 312 -19 709
rect 19 312 25 709
rect -25 300 25 312
rect -25 -312 25 -300
rect -25 -709 -19 -312
rect 19 -709 25 -312
rect -25 -721 25 -709
<< res0p35 >>
rect -37 -297 37 297
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string parameters w 0.350 l 2.95 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 2.805k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 0.350 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
