magic
tech sky130A
magscale 1 2
timestamp 1628068563
<< error_p >>
rect -269 501 -211 507
rect -77 501 -19 507
rect 115 501 173 507
rect 307 501 365 507
rect -269 467 -257 501
rect -77 467 -65 501
rect 115 467 127 501
rect 307 467 319 501
rect -269 461 -211 467
rect -77 461 -19 467
rect 115 461 173 467
rect 307 461 365 467
rect -365 -467 -307 -461
rect -173 -467 -115 -461
rect 19 -467 77 -461
rect 211 -467 269 -461
rect -365 -501 -353 -467
rect -173 -501 -161 -467
rect 19 -501 31 -467
rect 211 -501 223 -467
rect -365 -507 -307 -501
rect -173 -507 -115 -501
rect 19 -507 77 -501
rect 211 -507 269 -501
<< nwell >>
rect -551 -639 551 639
<< pmos >>
rect -351 -420 -321 420
rect -255 -420 -225 420
rect -159 -420 -129 420
rect -63 -420 -33 420
rect 33 -420 63 420
rect 129 -420 159 420
rect 225 -420 255 420
rect 321 -420 351 420
<< pdiff >>
rect -413 408 -351 420
rect -413 -408 -401 408
rect -367 -408 -351 408
rect -413 -420 -351 -408
rect -321 408 -255 420
rect -321 -408 -305 408
rect -271 -408 -255 408
rect -321 -420 -255 -408
rect -225 408 -159 420
rect -225 -408 -209 408
rect -175 -408 -159 408
rect -225 -420 -159 -408
rect -129 408 -63 420
rect -129 -408 -113 408
rect -79 -408 -63 408
rect -129 -420 -63 -408
rect -33 408 33 420
rect -33 -408 -17 408
rect 17 -408 33 408
rect -33 -420 33 -408
rect 63 408 129 420
rect 63 -408 79 408
rect 113 -408 129 408
rect 63 -420 129 -408
rect 159 408 225 420
rect 159 -408 175 408
rect 209 -408 225 408
rect 159 -420 225 -408
rect 255 408 321 420
rect 255 -408 271 408
rect 305 -408 321 408
rect 255 -420 321 -408
rect 351 408 413 420
rect 351 -408 367 408
rect 401 -408 413 408
rect 351 -420 413 -408
<< pdiffc >>
rect -401 -408 -367 408
rect -305 -408 -271 408
rect -209 -408 -175 408
rect -113 -408 -79 408
rect -17 -408 17 408
rect 79 -408 113 408
rect 175 -408 209 408
rect 271 -408 305 408
rect 367 -408 401 408
<< nsubdiff >>
rect -515 569 -419 603
rect 419 569 515 603
rect -515 507 -481 569
rect 481 507 515 569
rect -515 -569 -481 -507
rect 481 -569 515 -507
rect -515 -603 -419 -569
rect 419 -603 515 -569
<< nsubdiffcont >>
rect -419 569 419 603
rect -515 -507 -481 507
rect 481 -507 515 507
rect -419 -603 419 -569
<< poly >>
rect -273 501 -207 517
rect -273 467 -257 501
rect -223 467 -207 501
rect -273 451 -207 467
rect -81 501 -15 517
rect -81 467 -65 501
rect -31 467 -15 501
rect -81 451 -15 467
rect 111 501 177 517
rect 111 467 127 501
rect 161 467 177 501
rect 111 451 177 467
rect 303 501 369 517
rect 303 467 319 501
rect 353 467 369 501
rect 303 451 369 467
rect -351 420 -321 446
rect -255 420 -225 451
rect -159 420 -129 446
rect -63 420 -33 451
rect 33 420 63 446
rect 129 420 159 451
rect 225 420 255 446
rect 321 420 351 451
rect -351 -451 -321 -420
rect -255 -446 -225 -420
rect -159 -451 -129 -420
rect -63 -446 -33 -420
rect 33 -451 63 -420
rect 129 -446 159 -420
rect 225 -451 255 -420
rect 321 -446 351 -420
rect -369 -467 -303 -451
rect -369 -501 -353 -467
rect -319 -501 -303 -467
rect -369 -517 -303 -501
rect -177 -467 -111 -451
rect -177 -501 -161 -467
rect -127 -501 -111 -467
rect -177 -517 -111 -501
rect 15 -467 81 -451
rect 15 -501 31 -467
rect 65 -501 81 -467
rect 15 -517 81 -501
rect 207 -467 273 -451
rect 207 -501 223 -467
rect 257 -501 273 -467
rect 207 -517 273 -501
<< polycont >>
rect -257 467 -223 501
rect -65 467 -31 501
rect 127 467 161 501
rect 319 467 353 501
rect -353 -501 -319 -467
rect -161 -501 -127 -467
rect 31 -501 65 -467
rect 223 -501 257 -467
<< locali >>
rect -515 569 -419 603
rect 419 569 515 603
rect -515 507 -481 569
rect 481 507 515 569
rect -273 467 -257 501
rect -223 467 -207 501
rect -81 467 -65 501
rect -31 467 -15 501
rect 111 467 127 501
rect 161 467 177 501
rect 303 467 319 501
rect 353 467 369 501
rect -401 408 -367 424
rect -401 -424 -367 -408
rect -305 408 -271 424
rect -305 -424 -271 -408
rect -209 408 -175 424
rect -209 -424 -175 -408
rect -113 408 -79 424
rect -113 -424 -79 -408
rect -17 408 17 424
rect -17 -424 17 -408
rect 79 408 113 424
rect 79 -424 113 -408
rect 175 408 209 424
rect 175 -424 209 -408
rect 271 408 305 424
rect 271 -424 305 -408
rect 367 408 401 424
rect 367 -424 401 -408
rect -369 -501 -353 -467
rect -319 -501 -303 -467
rect -177 -501 -161 -467
rect -127 -501 -111 -467
rect 15 -501 31 -467
rect 65 -501 81 -467
rect 207 -501 223 -467
rect 257 -501 273 -467
rect -515 -569 -481 -507
rect 481 -569 515 -507
rect -515 -603 -419 -569
rect 419 -603 515 -569
<< viali >>
rect -257 467 -223 501
rect -65 467 -31 501
rect 127 467 161 501
rect 319 467 353 501
rect -401 -408 -367 408
rect -305 -408 -271 408
rect -209 -408 -175 408
rect -113 -408 -79 408
rect -17 -408 17 408
rect 79 -408 113 408
rect 175 -408 209 408
rect 271 -408 305 408
rect 367 -408 401 408
rect -353 -501 -319 -467
rect -161 -501 -127 -467
rect 31 -501 65 -467
rect 223 -501 257 -467
<< metal1 >>
rect -269 501 -211 507
rect -269 467 -257 501
rect -223 467 -211 501
rect -269 461 -211 467
rect -77 501 -19 507
rect -77 467 -65 501
rect -31 467 -19 501
rect -77 461 -19 467
rect 115 501 173 507
rect 115 467 127 501
rect 161 467 173 501
rect 115 461 173 467
rect 307 501 365 507
rect 307 467 319 501
rect 353 467 365 501
rect 307 461 365 467
rect -407 408 -361 420
rect -407 -408 -401 408
rect -367 -408 -361 408
rect -407 -420 -361 -408
rect -311 408 -265 420
rect -311 -408 -305 408
rect -271 -408 -265 408
rect -311 -420 -265 -408
rect -215 408 -169 420
rect -215 -408 -209 408
rect -175 -408 -169 408
rect -215 -420 -169 -408
rect -119 408 -73 420
rect -119 -408 -113 408
rect -79 -408 -73 408
rect -119 -420 -73 -408
rect -23 408 23 420
rect -23 -408 -17 408
rect 17 -408 23 408
rect -23 -420 23 -408
rect 73 408 119 420
rect 73 -408 79 408
rect 113 -408 119 408
rect 73 -420 119 -408
rect 169 408 215 420
rect 169 -408 175 408
rect 209 -408 215 408
rect 169 -420 215 -408
rect 265 408 311 420
rect 265 -408 271 408
rect 305 -408 311 408
rect 265 -420 311 -408
rect 361 408 407 420
rect 361 -408 367 408
rect 401 -408 407 408
rect 361 -420 407 -408
rect -365 -467 -307 -461
rect -365 -501 -353 -467
rect -319 -501 -307 -467
rect -365 -507 -307 -501
rect -173 -467 -115 -461
rect -173 -501 -161 -467
rect -127 -501 -115 -467
rect -173 -507 -115 -501
rect 19 -467 77 -461
rect 19 -501 31 -467
rect 65 -501 77 -467
rect 19 -507 77 -501
rect 211 -467 269 -461
rect 211 -501 223 -467
rect 257 -501 269 -467
rect 211 -507 269 -501
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -498 -586 498 586
string parameters w 4.2 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
