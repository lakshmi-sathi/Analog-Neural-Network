magic
tech sky130A
magscale 1 2
timestamp 1626798771
<< error_p >>
rect -989 799 -931 805
rect -797 799 -739 805
rect -605 799 -547 805
rect -413 799 -355 805
rect -221 799 -163 805
rect -29 799 29 805
rect 163 799 221 805
rect 355 799 413 805
rect 547 799 605 805
rect 739 799 797 805
rect 931 799 989 805
rect -989 765 -977 799
rect -797 765 -785 799
rect -605 765 -593 799
rect -413 765 -401 799
rect -221 765 -209 799
rect -29 765 -17 799
rect 163 765 175 799
rect 355 765 367 799
rect 547 765 559 799
rect 739 765 751 799
rect 931 765 943 799
rect -989 759 -931 765
rect -797 759 -739 765
rect -605 759 -547 765
rect -413 759 -355 765
rect -221 759 -163 765
rect -29 759 29 765
rect 163 759 221 765
rect 355 759 413 765
rect 547 759 605 765
rect 739 759 797 765
rect 931 759 989 765
rect -893 71 -835 77
rect -701 71 -643 77
rect -509 71 -451 77
rect -317 71 -259 77
rect -125 71 -67 77
rect 67 71 125 77
rect 259 71 317 77
rect 451 71 509 77
rect 643 71 701 77
rect 835 71 893 77
rect -893 37 -881 71
rect -701 37 -689 71
rect -509 37 -497 71
rect -317 37 -305 71
rect -125 37 -113 71
rect 67 37 79 71
rect 259 37 271 71
rect 451 37 463 71
rect 643 37 655 71
rect 835 37 847 71
rect -893 31 -835 37
rect -701 31 -643 37
rect -509 31 -451 37
rect -317 31 -259 37
rect -125 31 -67 37
rect 67 31 125 37
rect 259 31 317 37
rect 451 31 509 37
rect 643 31 701 37
rect 835 31 893 37
rect -893 -37 -835 -31
rect -701 -37 -643 -31
rect -509 -37 -451 -31
rect -317 -37 -259 -31
rect -125 -37 -67 -31
rect 67 -37 125 -31
rect 259 -37 317 -31
rect 451 -37 509 -31
rect 643 -37 701 -31
rect 835 -37 893 -31
rect -893 -71 -881 -37
rect -701 -71 -689 -37
rect -509 -71 -497 -37
rect -317 -71 -305 -37
rect -125 -71 -113 -37
rect 67 -71 79 -37
rect 259 -71 271 -37
rect 451 -71 463 -37
rect 643 -71 655 -37
rect 835 -71 847 -37
rect -893 -77 -835 -71
rect -701 -77 -643 -71
rect -509 -77 -451 -71
rect -317 -77 -259 -71
rect -125 -77 -67 -71
rect 67 -77 125 -71
rect 259 -77 317 -71
rect 451 -77 509 -71
rect 643 -77 701 -71
rect 835 -77 893 -71
rect -989 -765 -931 -759
rect -797 -765 -739 -759
rect -605 -765 -547 -759
rect -413 -765 -355 -759
rect -221 -765 -163 -759
rect -29 -765 29 -759
rect 163 -765 221 -759
rect 355 -765 413 -759
rect 547 -765 605 -759
rect 739 -765 797 -759
rect 931 -765 989 -759
rect -989 -799 -977 -765
rect -797 -799 -785 -765
rect -605 -799 -593 -765
rect -413 -799 -401 -765
rect -221 -799 -209 -765
rect -29 -799 -17 -765
rect 163 -799 175 -765
rect 355 -799 367 -765
rect 547 -799 559 -765
rect 739 -799 751 -765
rect 931 -799 943 -765
rect -989 -805 -931 -799
rect -797 -805 -739 -799
rect -605 -805 -547 -799
rect -413 -805 -355 -799
rect -221 -805 -163 -799
rect -29 -805 29 -799
rect 163 -805 221 -799
rect 355 -805 413 -799
rect 547 -805 605 -799
rect 739 -805 797 -799
rect 931 -805 989 -799
<< nwell >>
rect -1175 -937 1175 937
<< pmos >>
rect -975 118 -945 718
rect -879 118 -849 718
rect -783 118 -753 718
rect -687 118 -657 718
rect -591 118 -561 718
rect -495 118 -465 718
rect -399 118 -369 718
rect -303 118 -273 718
rect -207 118 -177 718
rect -111 118 -81 718
rect -15 118 15 718
rect 81 118 111 718
rect 177 118 207 718
rect 273 118 303 718
rect 369 118 399 718
rect 465 118 495 718
rect 561 118 591 718
rect 657 118 687 718
rect 753 118 783 718
rect 849 118 879 718
rect 945 118 975 718
rect -975 -718 -945 -118
rect -879 -718 -849 -118
rect -783 -718 -753 -118
rect -687 -718 -657 -118
rect -591 -718 -561 -118
rect -495 -718 -465 -118
rect -399 -718 -369 -118
rect -303 -718 -273 -118
rect -207 -718 -177 -118
rect -111 -718 -81 -118
rect -15 -718 15 -118
rect 81 -718 111 -118
rect 177 -718 207 -118
rect 273 -718 303 -118
rect 369 -718 399 -118
rect 465 -718 495 -118
rect 561 -718 591 -118
rect 657 -718 687 -118
rect 753 -718 783 -118
rect 849 -718 879 -118
rect 945 -718 975 -118
<< pdiff >>
rect -1037 706 -975 718
rect -1037 130 -1025 706
rect -991 130 -975 706
rect -1037 118 -975 130
rect -945 706 -879 718
rect -945 130 -929 706
rect -895 130 -879 706
rect -945 118 -879 130
rect -849 706 -783 718
rect -849 130 -833 706
rect -799 130 -783 706
rect -849 118 -783 130
rect -753 706 -687 718
rect -753 130 -737 706
rect -703 130 -687 706
rect -753 118 -687 130
rect -657 706 -591 718
rect -657 130 -641 706
rect -607 130 -591 706
rect -657 118 -591 130
rect -561 706 -495 718
rect -561 130 -545 706
rect -511 130 -495 706
rect -561 118 -495 130
rect -465 706 -399 718
rect -465 130 -449 706
rect -415 130 -399 706
rect -465 118 -399 130
rect -369 706 -303 718
rect -369 130 -353 706
rect -319 130 -303 706
rect -369 118 -303 130
rect -273 706 -207 718
rect -273 130 -257 706
rect -223 130 -207 706
rect -273 118 -207 130
rect -177 706 -111 718
rect -177 130 -161 706
rect -127 130 -111 706
rect -177 118 -111 130
rect -81 706 -15 718
rect -81 130 -65 706
rect -31 130 -15 706
rect -81 118 -15 130
rect 15 706 81 718
rect 15 130 31 706
rect 65 130 81 706
rect 15 118 81 130
rect 111 706 177 718
rect 111 130 127 706
rect 161 130 177 706
rect 111 118 177 130
rect 207 706 273 718
rect 207 130 223 706
rect 257 130 273 706
rect 207 118 273 130
rect 303 706 369 718
rect 303 130 319 706
rect 353 130 369 706
rect 303 118 369 130
rect 399 706 465 718
rect 399 130 415 706
rect 449 130 465 706
rect 399 118 465 130
rect 495 706 561 718
rect 495 130 511 706
rect 545 130 561 706
rect 495 118 561 130
rect 591 706 657 718
rect 591 130 607 706
rect 641 130 657 706
rect 591 118 657 130
rect 687 706 753 718
rect 687 130 703 706
rect 737 130 753 706
rect 687 118 753 130
rect 783 706 849 718
rect 783 130 799 706
rect 833 130 849 706
rect 783 118 849 130
rect 879 706 945 718
rect 879 130 895 706
rect 929 130 945 706
rect 879 118 945 130
rect 975 706 1037 718
rect 975 130 991 706
rect 1025 130 1037 706
rect 975 118 1037 130
rect -1037 -130 -975 -118
rect -1037 -706 -1025 -130
rect -991 -706 -975 -130
rect -1037 -718 -975 -706
rect -945 -130 -879 -118
rect -945 -706 -929 -130
rect -895 -706 -879 -130
rect -945 -718 -879 -706
rect -849 -130 -783 -118
rect -849 -706 -833 -130
rect -799 -706 -783 -130
rect -849 -718 -783 -706
rect -753 -130 -687 -118
rect -753 -706 -737 -130
rect -703 -706 -687 -130
rect -753 -718 -687 -706
rect -657 -130 -591 -118
rect -657 -706 -641 -130
rect -607 -706 -591 -130
rect -657 -718 -591 -706
rect -561 -130 -495 -118
rect -561 -706 -545 -130
rect -511 -706 -495 -130
rect -561 -718 -495 -706
rect -465 -130 -399 -118
rect -465 -706 -449 -130
rect -415 -706 -399 -130
rect -465 -718 -399 -706
rect -369 -130 -303 -118
rect -369 -706 -353 -130
rect -319 -706 -303 -130
rect -369 -718 -303 -706
rect -273 -130 -207 -118
rect -273 -706 -257 -130
rect -223 -706 -207 -130
rect -273 -718 -207 -706
rect -177 -130 -111 -118
rect -177 -706 -161 -130
rect -127 -706 -111 -130
rect -177 -718 -111 -706
rect -81 -130 -15 -118
rect -81 -706 -65 -130
rect -31 -706 -15 -130
rect -81 -718 -15 -706
rect 15 -130 81 -118
rect 15 -706 31 -130
rect 65 -706 81 -130
rect 15 -718 81 -706
rect 111 -130 177 -118
rect 111 -706 127 -130
rect 161 -706 177 -130
rect 111 -718 177 -706
rect 207 -130 273 -118
rect 207 -706 223 -130
rect 257 -706 273 -130
rect 207 -718 273 -706
rect 303 -130 369 -118
rect 303 -706 319 -130
rect 353 -706 369 -130
rect 303 -718 369 -706
rect 399 -130 465 -118
rect 399 -706 415 -130
rect 449 -706 465 -130
rect 399 -718 465 -706
rect 495 -130 561 -118
rect 495 -706 511 -130
rect 545 -706 561 -130
rect 495 -718 561 -706
rect 591 -130 657 -118
rect 591 -706 607 -130
rect 641 -706 657 -130
rect 591 -718 657 -706
rect 687 -130 753 -118
rect 687 -706 703 -130
rect 737 -706 753 -130
rect 687 -718 753 -706
rect 783 -130 849 -118
rect 783 -706 799 -130
rect 833 -706 849 -130
rect 783 -718 849 -706
rect 879 -130 945 -118
rect 879 -706 895 -130
rect 929 -706 945 -130
rect 879 -718 945 -706
rect 975 -130 1037 -118
rect 975 -706 991 -130
rect 1025 -706 1037 -130
rect 975 -718 1037 -706
<< pdiffc >>
rect -1025 130 -991 706
rect -929 130 -895 706
rect -833 130 -799 706
rect -737 130 -703 706
rect -641 130 -607 706
rect -545 130 -511 706
rect -449 130 -415 706
rect -353 130 -319 706
rect -257 130 -223 706
rect -161 130 -127 706
rect -65 130 -31 706
rect 31 130 65 706
rect 127 130 161 706
rect 223 130 257 706
rect 319 130 353 706
rect 415 130 449 706
rect 511 130 545 706
rect 607 130 641 706
rect 703 130 737 706
rect 799 130 833 706
rect 895 130 929 706
rect 991 130 1025 706
rect -1025 -706 -991 -130
rect -929 -706 -895 -130
rect -833 -706 -799 -130
rect -737 -706 -703 -130
rect -641 -706 -607 -130
rect -545 -706 -511 -130
rect -449 -706 -415 -130
rect -353 -706 -319 -130
rect -257 -706 -223 -130
rect -161 -706 -127 -130
rect -65 -706 -31 -130
rect 31 -706 65 -130
rect 127 -706 161 -130
rect 223 -706 257 -130
rect 319 -706 353 -130
rect 415 -706 449 -130
rect 511 -706 545 -130
rect 607 -706 641 -130
rect 703 -706 737 -130
rect 799 -706 833 -130
rect 895 -706 929 -130
rect 991 -706 1025 -130
<< nsubdiff >>
rect -1139 867 -1043 901
rect 1043 867 1139 901
rect -1139 805 -1105 867
rect 1105 805 1139 867
rect -1139 -867 -1105 -805
rect 1105 -867 1139 -805
rect -1139 -901 -1043 -867
rect 1043 -901 1139 -867
<< nsubdiffcont >>
rect -1043 867 1043 901
rect -1139 -805 -1105 805
rect 1105 -805 1139 805
rect -1043 -901 1043 -867
<< poly >>
rect -993 799 -927 815
rect -993 765 -977 799
rect -943 765 -927 799
rect -993 749 -927 765
rect -801 799 -735 815
rect -801 765 -785 799
rect -751 765 -735 799
rect -801 749 -735 765
rect -609 799 -543 815
rect -609 765 -593 799
rect -559 765 -543 799
rect -609 749 -543 765
rect -417 799 -351 815
rect -417 765 -401 799
rect -367 765 -351 799
rect -417 749 -351 765
rect -225 799 -159 815
rect -225 765 -209 799
rect -175 765 -159 799
rect -225 749 -159 765
rect -33 799 33 815
rect -33 765 -17 799
rect 17 765 33 799
rect -33 749 33 765
rect 159 799 225 815
rect 159 765 175 799
rect 209 765 225 799
rect 159 749 225 765
rect 351 799 417 815
rect 351 765 367 799
rect 401 765 417 799
rect 351 749 417 765
rect 543 799 609 815
rect 543 765 559 799
rect 593 765 609 799
rect 543 749 609 765
rect 735 799 801 815
rect 735 765 751 799
rect 785 765 801 799
rect 735 749 801 765
rect 927 799 993 815
rect 927 765 943 799
rect 977 765 993 799
rect 927 749 993 765
rect -975 718 -945 749
rect -879 718 -849 744
rect -783 718 -753 749
rect -687 718 -657 744
rect -591 718 -561 749
rect -495 718 -465 744
rect -399 718 -369 749
rect -303 718 -273 744
rect -207 718 -177 749
rect -111 718 -81 744
rect -15 718 15 749
rect 81 718 111 744
rect 177 718 207 749
rect 273 718 303 744
rect 369 718 399 749
rect 465 718 495 744
rect 561 718 591 749
rect 657 718 687 744
rect 753 718 783 749
rect 849 718 879 744
rect 945 718 975 749
rect -975 92 -945 118
rect -879 87 -849 118
rect -783 92 -753 118
rect -687 87 -657 118
rect -591 92 -561 118
rect -495 87 -465 118
rect -399 92 -369 118
rect -303 87 -273 118
rect -207 92 -177 118
rect -111 87 -81 118
rect -15 92 15 118
rect 81 87 111 118
rect 177 92 207 118
rect 273 87 303 118
rect 369 92 399 118
rect 465 87 495 118
rect 561 92 591 118
rect 657 87 687 118
rect 753 92 783 118
rect 849 87 879 118
rect 945 92 975 118
rect -897 71 -831 87
rect -897 37 -881 71
rect -847 37 -831 71
rect -897 21 -831 37
rect -705 71 -639 87
rect -705 37 -689 71
rect -655 37 -639 71
rect -705 21 -639 37
rect -513 71 -447 87
rect -513 37 -497 71
rect -463 37 -447 71
rect -513 21 -447 37
rect -321 71 -255 87
rect -321 37 -305 71
rect -271 37 -255 71
rect -321 21 -255 37
rect -129 71 -63 87
rect -129 37 -113 71
rect -79 37 -63 71
rect -129 21 -63 37
rect 63 71 129 87
rect 63 37 79 71
rect 113 37 129 71
rect 63 21 129 37
rect 255 71 321 87
rect 255 37 271 71
rect 305 37 321 71
rect 255 21 321 37
rect 447 71 513 87
rect 447 37 463 71
rect 497 37 513 71
rect 447 21 513 37
rect 639 71 705 87
rect 639 37 655 71
rect 689 37 705 71
rect 639 21 705 37
rect 831 71 897 87
rect 831 37 847 71
rect 881 37 897 71
rect 831 21 897 37
rect -897 -37 -831 -21
rect -897 -71 -881 -37
rect -847 -71 -831 -37
rect -897 -87 -831 -71
rect -705 -37 -639 -21
rect -705 -71 -689 -37
rect -655 -71 -639 -37
rect -705 -87 -639 -71
rect -513 -37 -447 -21
rect -513 -71 -497 -37
rect -463 -71 -447 -37
rect -513 -87 -447 -71
rect -321 -37 -255 -21
rect -321 -71 -305 -37
rect -271 -71 -255 -37
rect -321 -87 -255 -71
rect -129 -37 -63 -21
rect -129 -71 -113 -37
rect -79 -71 -63 -37
rect -129 -87 -63 -71
rect 63 -37 129 -21
rect 63 -71 79 -37
rect 113 -71 129 -37
rect 63 -87 129 -71
rect 255 -37 321 -21
rect 255 -71 271 -37
rect 305 -71 321 -37
rect 255 -87 321 -71
rect 447 -37 513 -21
rect 447 -71 463 -37
rect 497 -71 513 -37
rect 447 -87 513 -71
rect 639 -37 705 -21
rect 639 -71 655 -37
rect 689 -71 705 -37
rect 639 -87 705 -71
rect 831 -37 897 -21
rect 831 -71 847 -37
rect 881 -71 897 -37
rect 831 -87 897 -71
rect -975 -118 -945 -92
rect -879 -118 -849 -87
rect -783 -118 -753 -92
rect -687 -118 -657 -87
rect -591 -118 -561 -92
rect -495 -118 -465 -87
rect -399 -118 -369 -92
rect -303 -118 -273 -87
rect -207 -118 -177 -92
rect -111 -118 -81 -87
rect -15 -118 15 -92
rect 81 -118 111 -87
rect 177 -118 207 -92
rect 273 -118 303 -87
rect 369 -118 399 -92
rect 465 -118 495 -87
rect 561 -118 591 -92
rect 657 -118 687 -87
rect 753 -118 783 -92
rect 849 -118 879 -87
rect 945 -118 975 -92
rect -975 -749 -945 -718
rect -879 -744 -849 -718
rect -783 -749 -753 -718
rect -687 -744 -657 -718
rect -591 -749 -561 -718
rect -495 -744 -465 -718
rect -399 -749 -369 -718
rect -303 -744 -273 -718
rect -207 -749 -177 -718
rect -111 -744 -81 -718
rect -15 -749 15 -718
rect 81 -744 111 -718
rect 177 -749 207 -718
rect 273 -744 303 -718
rect 369 -749 399 -718
rect 465 -744 495 -718
rect 561 -749 591 -718
rect 657 -744 687 -718
rect 753 -749 783 -718
rect 849 -744 879 -718
rect 945 -749 975 -718
rect -993 -765 -927 -749
rect -993 -799 -977 -765
rect -943 -799 -927 -765
rect -993 -815 -927 -799
rect -801 -765 -735 -749
rect -801 -799 -785 -765
rect -751 -799 -735 -765
rect -801 -815 -735 -799
rect -609 -765 -543 -749
rect -609 -799 -593 -765
rect -559 -799 -543 -765
rect -609 -815 -543 -799
rect -417 -765 -351 -749
rect -417 -799 -401 -765
rect -367 -799 -351 -765
rect -417 -815 -351 -799
rect -225 -765 -159 -749
rect -225 -799 -209 -765
rect -175 -799 -159 -765
rect -225 -815 -159 -799
rect -33 -765 33 -749
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -815 33 -799
rect 159 -765 225 -749
rect 159 -799 175 -765
rect 209 -799 225 -765
rect 159 -815 225 -799
rect 351 -765 417 -749
rect 351 -799 367 -765
rect 401 -799 417 -765
rect 351 -815 417 -799
rect 543 -765 609 -749
rect 543 -799 559 -765
rect 593 -799 609 -765
rect 543 -815 609 -799
rect 735 -765 801 -749
rect 735 -799 751 -765
rect 785 -799 801 -765
rect 735 -815 801 -799
rect 927 -765 993 -749
rect 927 -799 943 -765
rect 977 -799 993 -765
rect 927 -815 993 -799
<< polycont >>
rect -977 765 -943 799
rect -785 765 -751 799
rect -593 765 -559 799
rect -401 765 -367 799
rect -209 765 -175 799
rect -17 765 17 799
rect 175 765 209 799
rect 367 765 401 799
rect 559 765 593 799
rect 751 765 785 799
rect 943 765 977 799
rect -881 37 -847 71
rect -689 37 -655 71
rect -497 37 -463 71
rect -305 37 -271 71
rect -113 37 -79 71
rect 79 37 113 71
rect 271 37 305 71
rect 463 37 497 71
rect 655 37 689 71
rect 847 37 881 71
rect -881 -71 -847 -37
rect -689 -71 -655 -37
rect -497 -71 -463 -37
rect -305 -71 -271 -37
rect -113 -71 -79 -37
rect 79 -71 113 -37
rect 271 -71 305 -37
rect 463 -71 497 -37
rect 655 -71 689 -37
rect 847 -71 881 -37
rect -977 -799 -943 -765
rect -785 -799 -751 -765
rect -593 -799 -559 -765
rect -401 -799 -367 -765
rect -209 -799 -175 -765
rect -17 -799 17 -765
rect 175 -799 209 -765
rect 367 -799 401 -765
rect 559 -799 593 -765
rect 751 -799 785 -765
rect 943 -799 977 -765
<< locali >>
rect -1139 867 -1043 901
rect 1043 867 1139 901
rect -1139 805 -1105 867
rect 1105 805 1139 867
rect -993 765 -977 799
rect -943 765 -927 799
rect -801 765 -785 799
rect -751 765 -735 799
rect -609 765 -593 799
rect -559 765 -543 799
rect -417 765 -401 799
rect -367 765 -351 799
rect -225 765 -209 799
rect -175 765 -159 799
rect -33 765 -17 799
rect 17 765 33 799
rect 159 765 175 799
rect 209 765 225 799
rect 351 765 367 799
rect 401 765 417 799
rect 543 765 559 799
rect 593 765 609 799
rect 735 765 751 799
rect 785 765 801 799
rect 927 765 943 799
rect 977 765 993 799
rect -1025 706 -991 722
rect -1025 114 -991 130
rect -929 706 -895 722
rect -929 114 -895 130
rect -833 706 -799 722
rect -833 114 -799 130
rect -737 706 -703 722
rect -737 114 -703 130
rect -641 706 -607 722
rect -641 114 -607 130
rect -545 706 -511 722
rect -545 114 -511 130
rect -449 706 -415 722
rect -449 114 -415 130
rect -353 706 -319 722
rect -353 114 -319 130
rect -257 706 -223 722
rect -257 114 -223 130
rect -161 706 -127 722
rect -161 114 -127 130
rect -65 706 -31 722
rect -65 114 -31 130
rect 31 706 65 722
rect 31 114 65 130
rect 127 706 161 722
rect 127 114 161 130
rect 223 706 257 722
rect 223 114 257 130
rect 319 706 353 722
rect 319 114 353 130
rect 415 706 449 722
rect 415 114 449 130
rect 511 706 545 722
rect 511 114 545 130
rect 607 706 641 722
rect 607 114 641 130
rect 703 706 737 722
rect 703 114 737 130
rect 799 706 833 722
rect 799 114 833 130
rect 895 706 929 722
rect 895 114 929 130
rect 991 706 1025 722
rect 991 114 1025 130
rect -897 37 -881 71
rect -847 37 -831 71
rect -705 37 -689 71
rect -655 37 -639 71
rect -513 37 -497 71
rect -463 37 -447 71
rect -321 37 -305 71
rect -271 37 -255 71
rect -129 37 -113 71
rect -79 37 -63 71
rect 63 37 79 71
rect 113 37 129 71
rect 255 37 271 71
rect 305 37 321 71
rect 447 37 463 71
rect 497 37 513 71
rect 639 37 655 71
rect 689 37 705 71
rect 831 37 847 71
rect 881 37 897 71
rect -897 -71 -881 -37
rect -847 -71 -831 -37
rect -705 -71 -689 -37
rect -655 -71 -639 -37
rect -513 -71 -497 -37
rect -463 -71 -447 -37
rect -321 -71 -305 -37
rect -271 -71 -255 -37
rect -129 -71 -113 -37
rect -79 -71 -63 -37
rect 63 -71 79 -37
rect 113 -71 129 -37
rect 255 -71 271 -37
rect 305 -71 321 -37
rect 447 -71 463 -37
rect 497 -71 513 -37
rect 639 -71 655 -37
rect 689 -71 705 -37
rect 831 -71 847 -37
rect 881 -71 897 -37
rect -1025 -130 -991 -114
rect -1025 -722 -991 -706
rect -929 -130 -895 -114
rect -929 -722 -895 -706
rect -833 -130 -799 -114
rect -833 -722 -799 -706
rect -737 -130 -703 -114
rect -737 -722 -703 -706
rect -641 -130 -607 -114
rect -641 -722 -607 -706
rect -545 -130 -511 -114
rect -545 -722 -511 -706
rect -449 -130 -415 -114
rect -449 -722 -415 -706
rect -353 -130 -319 -114
rect -353 -722 -319 -706
rect -257 -130 -223 -114
rect -257 -722 -223 -706
rect -161 -130 -127 -114
rect -161 -722 -127 -706
rect -65 -130 -31 -114
rect -65 -722 -31 -706
rect 31 -130 65 -114
rect 31 -722 65 -706
rect 127 -130 161 -114
rect 127 -722 161 -706
rect 223 -130 257 -114
rect 223 -722 257 -706
rect 319 -130 353 -114
rect 319 -722 353 -706
rect 415 -130 449 -114
rect 415 -722 449 -706
rect 511 -130 545 -114
rect 511 -722 545 -706
rect 607 -130 641 -114
rect 607 -722 641 -706
rect 703 -130 737 -114
rect 703 -722 737 -706
rect 799 -130 833 -114
rect 799 -722 833 -706
rect 895 -130 929 -114
rect 895 -722 929 -706
rect 991 -130 1025 -114
rect 991 -722 1025 -706
rect -993 -799 -977 -765
rect -943 -799 -927 -765
rect -801 -799 -785 -765
rect -751 -799 -735 -765
rect -609 -799 -593 -765
rect -559 -799 -543 -765
rect -417 -799 -401 -765
rect -367 -799 -351 -765
rect -225 -799 -209 -765
rect -175 -799 -159 -765
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect 159 -799 175 -765
rect 209 -799 225 -765
rect 351 -799 367 -765
rect 401 -799 417 -765
rect 543 -799 559 -765
rect 593 -799 609 -765
rect 735 -799 751 -765
rect 785 -799 801 -765
rect 927 -799 943 -765
rect 977 -799 993 -765
rect -1139 -867 -1105 -805
rect 1105 -867 1139 -805
rect -1139 -901 -1043 -867
rect 1043 -901 1139 -867
<< viali >>
rect -977 765 -943 799
rect -785 765 -751 799
rect -593 765 -559 799
rect -401 765 -367 799
rect -209 765 -175 799
rect -17 765 17 799
rect 175 765 209 799
rect 367 765 401 799
rect 559 765 593 799
rect 751 765 785 799
rect 943 765 977 799
rect -1025 130 -991 706
rect -929 130 -895 706
rect -833 130 -799 706
rect -737 130 -703 706
rect -641 130 -607 706
rect -545 130 -511 706
rect -449 130 -415 706
rect -353 130 -319 706
rect -257 130 -223 706
rect -161 130 -127 706
rect -65 130 -31 706
rect 31 130 65 706
rect 127 130 161 706
rect 223 130 257 706
rect 319 130 353 706
rect 415 130 449 706
rect 511 130 545 706
rect 607 130 641 706
rect 703 130 737 706
rect 799 130 833 706
rect 895 130 929 706
rect 991 130 1025 706
rect -881 37 -847 71
rect -689 37 -655 71
rect -497 37 -463 71
rect -305 37 -271 71
rect -113 37 -79 71
rect 79 37 113 71
rect 271 37 305 71
rect 463 37 497 71
rect 655 37 689 71
rect 847 37 881 71
rect -881 -71 -847 -37
rect -689 -71 -655 -37
rect -497 -71 -463 -37
rect -305 -71 -271 -37
rect -113 -71 -79 -37
rect 79 -71 113 -37
rect 271 -71 305 -37
rect 463 -71 497 -37
rect 655 -71 689 -37
rect 847 -71 881 -37
rect -1025 -706 -991 -130
rect -929 -706 -895 -130
rect -833 -706 -799 -130
rect -737 -706 -703 -130
rect -641 -706 -607 -130
rect -545 -706 -511 -130
rect -449 -706 -415 -130
rect -353 -706 -319 -130
rect -257 -706 -223 -130
rect -161 -706 -127 -130
rect -65 -706 -31 -130
rect 31 -706 65 -130
rect 127 -706 161 -130
rect 223 -706 257 -130
rect 319 -706 353 -130
rect 415 -706 449 -130
rect 511 -706 545 -130
rect 607 -706 641 -130
rect 703 -706 737 -130
rect 799 -706 833 -130
rect 895 -706 929 -130
rect 991 -706 1025 -130
rect -977 -799 -943 -765
rect -785 -799 -751 -765
rect -593 -799 -559 -765
rect -401 -799 -367 -765
rect -209 -799 -175 -765
rect -17 -799 17 -765
rect 175 -799 209 -765
rect 367 -799 401 -765
rect 559 -799 593 -765
rect 751 -799 785 -765
rect 943 -799 977 -765
<< metal1 >>
rect -989 799 -931 805
rect -989 765 -977 799
rect -943 765 -931 799
rect -989 759 -931 765
rect -797 799 -739 805
rect -797 765 -785 799
rect -751 765 -739 799
rect -797 759 -739 765
rect -605 799 -547 805
rect -605 765 -593 799
rect -559 765 -547 799
rect -605 759 -547 765
rect -413 799 -355 805
rect -413 765 -401 799
rect -367 765 -355 799
rect -413 759 -355 765
rect -221 799 -163 805
rect -221 765 -209 799
rect -175 765 -163 799
rect -221 759 -163 765
rect -29 799 29 805
rect -29 765 -17 799
rect 17 765 29 799
rect -29 759 29 765
rect 163 799 221 805
rect 163 765 175 799
rect 209 765 221 799
rect 163 759 221 765
rect 355 799 413 805
rect 355 765 367 799
rect 401 765 413 799
rect 355 759 413 765
rect 547 799 605 805
rect 547 765 559 799
rect 593 765 605 799
rect 547 759 605 765
rect 739 799 797 805
rect 739 765 751 799
rect 785 765 797 799
rect 739 759 797 765
rect 931 799 989 805
rect 931 765 943 799
rect 977 765 989 799
rect 931 759 989 765
rect -1031 706 -985 718
rect -1031 130 -1025 706
rect -991 130 -985 706
rect -1031 118 -985 130
rect -935 706 -889 718
rect -935 130 -929 706
rect -895 130 -889 706
rect -935 118 -889 130
rect -839 706 -793 718
rect -839 130 -833 706
rect -799 130 -793 706
rect -839 118 -793 130
rect -743 706 -697 718
rect -743 130 -737 706
rect -703 130 -697 706
rect -743 118 -697 130
rect -647 706 -601 718
rect -647 130 -641 706
rect -607 130 -601 706
rect -647 118 -601 130
rect -551 706 -505 718
rect -551 130 -545 706
rect -511 130 -505 706
rect -551 118 -505 130
rect -455 706 -409 718
rect -455 130 -449 706
rect -415 130 -409 706
rect -455 118 -409 130
rect -359 706 -313 718
rect -359 130 -353 706
rect -319 130 -313 706
rect -359 118 -313 130
rect -263 706 -217 718
rect -263 130 -257 706
rect -223 130 -217 706
rect -263 118 -217 130
rect -167 706 -121 718
rect -167 130 -161 706
rect -127 130 -121 706
rect -167 118 -121 130
rect -71 706 -25 718
rect -71 130 -65 706
rect -31 130 -25 706
rect -71 118 -25 130
rect 25 706 71 718
rect 25 130 31 706
rect 65 130 71 706
rect 25 118 71 130
rect 121 706 167 718
rect 121 130 127 706
rect 161 130 167 706
rect 121 118 167 130
rect 217 706 263 718
rect 217 130 223 706
rect 257 130 263 706
rect 217 118 263 130
rect 313 706 359 718
rect 313 130 319 706
rect 353 130 359 706
rect 313 118 359 130
rect 409 706 455 718
rect 409 130 415 706
rect 449 130 455 706
rect 409 118 455 130
rect 505 706 551 718
rect 505 130 511 706
rect 545 130 551 706
rect 505 118 551 130
rect 601 706 647 718
rect 601 130 607 706
rect 641 130 647 706
rect 601 118 647 130
rect 697 706 743 718
rect 697 130 703 706
rect 737 130 743 706
rect 697 118 743 130
rect 793 706 839 718
rect 793 130 799 706
rect 833 130 839 706
rect 793 118 839 130
rect 889 706 935 718
rect 889 130 895 706
rect 929 130 935 706
rect 889 118 935 130
rect 985 706 1031 718
rect 985 130 991 706
rect 1025 130 1031 706
rect 985 118 1031 130
rect -893 71 -835 77
rect -893 37 -881 71
rect -847 37 -835 71
rect -893 31 -835 37
rect -701 71 -643 77
rect -701 37 -689 71
rect -655 37 -643 71
rect -701 31 -643 37
rect -509 71 -451 77
rect -509 37 -497 71
rect -463 37 -451 71
rect -509 31 -451 37
rect -317 71 -259 77
rect -317 37 -305 71
rect -271 37 -259 71
rect -317 31 -259 37
rect -125 71 -67 77
rect -125 37 -113 71
rect -79 37 -67 71
rect -125 31 -67 37
rect 67 71 125 77
rect 67 37 79 71
rect 113 37 125 71
rect 67 31 125 37
rect 259 71 317 77
rect 259 37 271 71
rect 305 37 317 71
rect 259 31 317 37
rect 451 71 509 77
rect 451 37 463 71
rect 497 37 509 71
rect 451 31 509 37
rect 643 71 701 77
rect 643 37 655 71
rect 689 37 701 71
rect 643 31 701 37
rect 835 71 893 77
rect 835 37 847 71
rect 881 37 893 71
rect 835 31 893 37
rect -893 -37 -835 -31
rect -893 -71 -881 -37
rect -847 -71 -835 -37
rect -893 -77 -835 -71
rect -701 -37 -643 -31
rect -701 -71 -689 -37
rect -655 -71 -643 -37
rect -701 -77 -643 -71
rect -509 -37 -451 -31
rect -509 -71 -497 -37
rect -463 -71 -451 -37
rect -509 -77 -451 -71
rect -317 -37 -259 -31
rect -317 -71 -305 -37
rect -271 -71 -259 -37
rect -317 -77 -259 -71
rect -125 -37 -67 -31
rect -125 -71 -113 -37
rect -79 -71 -67 -37
rect -125 -77 -67 -71
rect 67 -37 125 -31
rect 67 -71 79 -37
rect 113 -71 125 -37
rect 67 -77 125 -71
rect 259 -37 317 -31
rect 259 -71 271 -37
rect 305 -71 317 -37
rect 259 -77 317 -71
rect 451 -37 509 -31
rect 451 -71 463 -37
rect 497 -71 509 -37
rect 451 -77 509 -71
rect 643 -37 701 -31
rect 643 -71 655 -37
rect 689 -71 701 -37
rect 643 -77 701 -71
rect 835 -37 893 -31
rect 835 -71 847 -37
rect 881 -71 893 -37
rect 835 -77 893 -71
rect -1031 -130 -985 -118
rect -1031 -706 -1025 -130
rect -991 -706 -985 -130
rect -1031 -718 -985 -706
rect -935 -130 -889 -118
rect -935 -706 -929 -130
rect -895 -706 -889 -130
rect -935 -718 -889 -706
rect -839 -130 -793 -118
rect -839 -706 -833 -130
rect -799 -706 -793 -130
rect -839 -718 -793 -706
rect -743 -130 -697 -118
rect -743 -706 -737 -130
rect -703 -706 -697 -130
rect -743 -718 -697 -706
rect -647 -130 -601 -118
rect -647 -706 -641 -130
rect -607 -706 -601 -130
rect -647 -718 -601 -706
rect -551 -130 -505 -118
rect -551 -706 -545 -130
rect -511 -706 -505 -130
rect -551 -718 -505 -706
rect -455 -130 -409 -118
rect -455 -706 -449 -130
rect -415 -706 -409 -130
rect -455 -718 -409 -706
rect -359 -130 -313 -118
rect -359 -706 -353 -130
rect -319 -706 -313 -130
rect -359 -718 -313 -706
rect -263 -130 -217 -118
rect -263 -706 -257 -130
rect -223 -706 -217 -130
rect -263 -718 -217 -706
rect -167 -130 -121 -118
rect -167 -706 -161 -130
rect -127 -706 -121 -130
rect -167 -718 -121 -706
rect -71 -130 -25 -118
rect -71 -706 -65 -130
rect -31 -706 -25 -130
rect -71 -718 -25 -706
rect 25 -130 71 -118
rect 25 -706 31 -130
rect 65 -706 71 -130
rect 25 -718 71 -706
rect 121 -130 167 -118
rect 121 -706 127 -130
rect 161 -706 167 -130
rect 121 -718 167 -706
rect 217 -130 263 -118
rect 217 -706 223 -130
rect 257 -706 263 -130
rect 217 -718 263 -706
rect 313 -130 359 -118
rect 313 -706 319 -130
rect 353 -706 359 -130
rect 313 -718 359 -706
rect 409 -130 455 -118
rect 409 -706 415 -130
rect 449 -706 455 -130
rect 409 -718 455 -706
rect 505 -130 551 -118
rect 505 -706 511 -130
rect 545 -706 551 -130
rect 505 -718 551 -706
rect 601 -130 647 -118
rect 601 -706 607 -130
rect 641 -706 647 -130
rect 601 -718 647 -706
rect 697 -130 743 -118
rect 697 -706 703 -130
rect 737 -706 743 -130
rect 697 -718 743 -706
rect 793 -130 839 -118
rect 793 -706 799 -130
rect 833 -706 839 -130
rect 793 -718 839 -706
rect 889 -130 935 -118
rect 889 -706 895 -130
rect 929 -706 935 -130
rect 889 -718 935 -706
rect 985 -130 1031 -118
rect 985 -706 991 -130
rect 1025 -706 1031 -130
rect 985 -718 1031 -706
rect -989 -765 -931 -759
rect -989 -799 -977 -765
rect -943 -799 -931 -765
rect -989 -805 -931 -799
rect -797 -765 -739 -759
rect -797 -799 -785 -765
rect -751 -799 -739 -765
rect -797 -805 -739 -799
rect -605 -765 -547 -759
rect -605 -799 -593 -765
rect -559 -799 -547 -765
rect -605 -805 -547 -799
rect -413 -765 -355 -759
rect -413 -799 -401 -765
rect -367 -799 -355 -765
rect -413 -805 -355 -799
rect -221 -765 -163 -759
rect -221 -799 -209 -765
rect -175 -799 -163 -765
rect -221 -805 -163 -799
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -805 29 -799
rect 163 -765 221 -759
rect 163 -799 175 -765
rect 209 -799 221 -765
rect 163 -805 221 -799
rect 355 -765 413 -759
rect 355 -799 367 -765
rect 401 -799 413 -765
rect 355 -805 413 -799
rect 547 -765 605 -759
rect 547 -799 559 -765
rect 593 -799 605 -765
rect 547 -805 605 -799
rect 739 -765 797 -759
rect 739 -799 751 -765
rect 785 -799 797 -765
rect 739 -805 797 -799
rect 931 -765 989 -759
rect 931 -799 943 -765
rect 977 -799 989 -765
rect 931 -805 989 -799
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1122 -884 1122 884
string parameters w 3 l 0.15 m 2 nf 21 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
