magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 343 35 775
rect -35 -775 35 -343
<< xpolyres >>
rect -35 -343 35 343
<< viali >>
rect -17 721 17 755
rect -17 649 17 683
rect -17 577 17 611
rect -17 505 17 539
rect -17 433 17 467
rect -17 361 17 395
rect -17 -396 17 -362
rect -17 -468 17 -434
rect -17 -540 17 -506
rect -17 -612 17 -578
rect -17 -684 17 -650
rect -17 -756 17 -722
<< metal1 >>
rect -25 755 25 769
rect -25 721 -17 755
rect 17 721 25 755
rect -25 683 25 721
rect -25 649 -17 683
rect 17 649 25 683
rect -25 611 25 649
rect -25 577 -17 611
rect 17 577 25 611
rect -25 539 25 577
rect -25 505 -17 539
rect 17 505 25 539
rect -25 467 25 505
rect -25 433 -17 467
rect 17 433 25 467
rect -25 395 25 433
rect -25 361 -17 395
rect 17 361 25 395
rect -25 348 25 361
rect -25 -362 25 -348
rect -25 -396 -17 -362
rect 17 -396 25 -362
rect -25 -434 25 -396
rect -25 -468 -17 -434
rect 17 -468 25 -434
rect -25 -506 25 -468
rect -25 -540 -17 -506
rect 17 -540 25 -506
rect -25 -578 25 -540
rect -25 -612 -17 -578
rect 17 -612 25 -578
rect -25 -650 25 -612
rect -25 -684 -17 -650
rect 17 -684 25 -650
rect -25 -722 25 -684
rect -25 -756 -17 -722
rect 17 -756 25 -722
rect -25 -769 25 -756
<< end >>
