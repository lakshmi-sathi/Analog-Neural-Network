magic
tech sky130A
magscale 1 2
timestamp 1628056522
<< error_p >>
rect -29 881 29 887
rect -29 847 -17 881
rect -29 841 29 847
<< pwell >>
rect -211 -1019 211 1019
<< nmos >>
rect -15 -871 15 809
<< ndiff >>
rect -73 797 -15 809
rect -73 -859 -61 797
rect -27 -859 -15 797
rect -73 -871 -15 -859
rect 15 797 73 809
rect 15 -859 27 797
rect 61 -859 73 797
rect 15 -871 73 -859
<< ndiffc >>
rect -61 -859 -27 797
rect 27 -859 61 797
<< psubdiff >>
rect -175 949 -79 983
rect 79 949 175 983
rect -175 887 -141 949
rect 141 887 175 949
rect -175 -949 -141 -887
rect 141 -949 175 -887
rect -175 -983 -79 -949
rect 79 -983 175 -949
<< psubdiffcont >>
rect -79 949 79 983
rect -175 -887 -141 887
rect 141 -887 175 887
rect -79 -983 79 -949
<< poly >>
rect -33 881 33 897
rect -33 847 -17 881
rect 17 847 33 881
rect -33 831 33 847
rect -15 809 15 831
rect -15 -897 15 -871
<< polycont >>
rect -17 847 17 881
<< locali >>
rect -175 949 -79 983
rect 79 949 175 983
rect -175 887 -141 949
rect 141 887 175 949
rect -33 847 -17 881
rect 17 847 33 881
rect -61 797 -27 813
rect -61 -875 -27 -859
rect 27 797 61 813
rect 27 -875 61 -859
rect -175 -949 -141 -887
rect 141 -949 175 -887
rect -175 -983 -79 -949
rect 79 -983 175 -949
<< viali >>
rect -17 847 17 881
rect -61 -859 -27 797
rect 27 -859 61 797
<< metal1 >>
rect -29 881 29 887
rect -29 847 -17 881
rect 17 847 29 881
rect -29 841 29 847
rect -67 797 -21 809
rect -67 -859 -61 797
rect -27 -859 -21 797
rect -67 -871 -21 -859
rect 21 797 67 809
rect 21 -859 27 797
rect 61 -859 67 797
rect 21 -871 67 -859
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -966 158 966
string parameters w 8.4 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
