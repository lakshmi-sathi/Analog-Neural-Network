magic
tech sky130A
magscale 1 2
timestamp 1627900655
<< metal1 >>
rect 34 7678 44 8190
rect 454 7678 464 8190
rect 34608 7624 34618 8322
rect 35182 7624 35192 8322
rect 68926 8282 69410 8292
rect 68926 7730 68962 8282
rect 69396 7730 69410 8282
rect 68926 7664 69410 7730
rect 18 4240 28 4726
rect 444 4240 454 4726
rect 34714 4230 34724 4734
rect 35122 4230 35132 4734
rect 68966 4250 68976 4738
rect 69414 4250 69424 4738
rect 32527 1952 35228 1958
rect 28 1452 38 1930
rect 470 1452 480 1930
rect 32527 1424 32552 1952
rect 32992 1424 35228 1952
rect 32527 1416 35228 1424
rect 66955 1918 69781 1962
rect 66955 1476 67046 1918
rect 67496 1476 69781 1918
rect 66955 1420 69781 1476
rect 32513 -1474 35230 -1463
rect 46 -1986 56 -1484
rect 504 -1986 514 -1484
rect 32513 -2002 32570 -1474
rect 33010 -2002 35230 -1474
rect 68976 -1972 68986 -1496
rect 69404 -1972 69414 -1496
rect 32513 -2005 35230 -2002
rect 20 -4796 30 -4324
rect 440 -4796 450 -4324
rect 34726 -4796 34736 -4302
rect 35036 -4796 35046 -4302
rect 68976 -4784 68986 -4296
rect 69424 -4784 69434 -4296
rect 66961 -7724 69573 -7709
rect 72 -8234 82 -7728
rect 432 -8234 442 -7728
rect 34730 -8240 34740 -7758
rect 35126 -8240 35136 -7758
rect 66961 -8242 66992 -7724
rect 67518 -8242 69573 -7724
rect 66961 -8251 69573 -8242
rect -32 -11212 -22 -10754
rect 344 -11212 354 -10754
rect 34642 -11260 34652 -10764
rect 35046 -11260 35056 -10764
rect -58 -14682 -48 -14180
rect 294 -14682 304 -14180
rect 34632 -14672 34642 -14192
rect 35026 -14672 35036 -14192
rect -80 -17496 -70 -16974
rect 310 -17496 320 -16974
rect 34598 -17502 34608 -16998
rect 35046 -17502 35056 -16998
<< via1 >>
rect 44 7678 454 8190
rect 34618 7624 35182 8322
rect 68962 7730 69396 8282
rect 28 4240 444 4726
rect 34724 4230 35122 4734
rect 68976 4250 69414 4738
rect 38 1452 470 1930
rect 32552 1424 32992 1952
rect 67046 1476 67496 1918
rect 56 -1986 504 -1484
rect 32570 -2002 33010 -1474
rect 68986 -1972 69404 -1496
rect 30 -4796 440 -4324
rect 34736 -4796 35036 -4302
rect 68986 -4784 69424 -4296
rect 82 -8234 432 -7728
rect 34740 -8240 35126 -7758
rect 66992 -8242 67518 -7724
rect -22 -11212 344 -10754
rect 34652 -11260 35046 -10764
rect -48 -14682 294 -14180
rect 34642 -14672 35026 -14192
rect -70 -17496 310 -16974
rect 34608 -17502 35046 -16998
<< metal2 >>
rect 1460 9280 99566 9417
rect 34618 8322 35182 8332
rect 44 8190 454 8200
rect 44 7668 454 7678
rect 68962 8282 69396 8292
rect 68962 7720 69396 7730
rect 34618 7614 35182 7624
rect 64882 5866 65228 5876
rect 30222 5844 30564 5854
rect 30222 5540 30564 5550
rect 64882 5540 65228 5550
rect 28 4726 444 4736
rect 28 4230 444 4240
rect 34724 4734 35122 4744
rect 68976 4738 69414 4748
rect 68976 4240 69414 4250
rect 34724 4220 35122 4230
rect -8550 1458 -7096 2048
rect -5372 1938 -4186 1953
rect 32552 1952 32992 1962
rect 38 1938 470 1940
rect -5382 1930 470 1938
rect -5382 1480 38 1930
rect -8550 -100 -8362 1458
rect -7296 -100 -7096 1458
rect -8550 -546 -7096 -100
rect -5372 -1484 -4186 1480
rect 38 1442 470 1452
rect 67046 1918 67496 1928
rect 67046 1466 67496 1476
rect 32552 1414 32992 1424
rect 28944 238 28966 240
rect 28944 120 28974 238
rect 2022 56 19190 110
rect 2022 -150 13690 56
rect 14226 -150 19190 56
rect 21204 94 28986 120
rect 63638 100 63664 294
rect 97884 124 97912 242
rect 21204 -26 54118 94
rect 21204 -140 48476 -26
rect 28658 -156 48476 -140
rect 13690 -212 14226 -202
rect 28944 -268 28974 -156
rect 28946 -274 28974 -268
rect 48456 -266 48476 -156
rect 48970 -156 54118 -26
rect 48970 -266 48992 -156
rect 55562 -162 88342 100
rect 48456 -288 48992 -266
rect 63638 -276 63664 -162
rect 89808 -170 97912 124
rect 97884 -282 97912 -170
rect 32570 -1474 33010 -1464
rect 56 -1484 504 -1474
rect -5372 -1958 56 -1484
rect -8612 -5478 -7158 -4846
rect -8612 -6996 -8406 -5478
rect -7286 -6996 -7158 -5478
rect -8612 -7440 -7158 -6996
rect -8550 -11908 -7096 -11172
rect -5372 -11908 -4186 -1958
rect 56 -1996 504 -1986
rect 68986 -1496 69404 -1486
rect 68986 -1982 69404 -1972
rect 32570 -2012 33010 -2002
rect 34736 -4302 35036 -4292
rect 30 -4324 440 -4314
rect 30 -4806 440 -4796
rect 68986 -4296 69424 -4286
rect 68986 -4794 69424 -4784
rect 34736 -4806 35036 -4796
rect 30208 -5580 30568 -5570
rect 30208 -5906 30568 -5896
rect 64870 -5584 65252 -5574
rect 64870 -6034 65252 -6024
rect 99112 -6733 99518 6411
rect 82 -7728 432 -7718
rect 66992 -7724 67518 -7714
rect 82 -8244 432 -8234
rect 34740 -7758 35126 -7748
rect 34740 -8250 35126 -8240
rect 66992 -8252 67518 -8242
rect 644 -9344 1786 -9338
rect 644 -9604 1778 -9344
rect 4370 -9378 30488 -9338
rect 4370 -9600 36660 -9378
rect 4362 -9604 36660 -9600
rect 28836 -9628 36660 -9604
rect 38876 -9628 99490 -9378
rect -22 -10754 344 -10744
rect -22 -11222 344 -11212
rect 34652 -10764 35046 -10754
rect 34652 -11270 35046 -11260
rect -8550 -13094 -4186 -11908
rect -8550 -13126 -6654 -13094
rect -8550 -13766 -7096 -13126
rect -5372 -16978 -4186 -13094
rect -48 -14180 294 -14170
rect 34642 -14192 35026 -14182
rect 34642 -14682 35026 -14672
rect -48 -14692 294 -14682
rect -70 -16974 310 -16964
rect -5372 -17476 -70 -16978
rect -5372 -17661 -4186 -17476
rect -70 -17506 310 -17496
rect 34608 -16998 35046 -16988
rect 34608 -17512 35046 -17502
rect 48434 -18612 49004 -18582
rect 13674 -18696 14250 -18686
rect 2038 -18910 13674 -18808
rect 48434 -18808 48494 -18612
rect 14250 -18870 48494 -18808
rect 48944 -18808 49004 -18612
rect 48944 -18870 63550 -18808
rect 14250 -18910 63550 -18870
rect 2038 -18920 63550 -18910
<< via2 >>
rect 44 7678 454 8190
rect 34618 7624 35182 8322
rect 68962 7730 69396 8282
rect 30222 5550 30564 5844
rect 64882 5550 65228 5866
rect 28 4240 444 4726
rect 34724 4230 35122 4734
rect 68976 4250 69414 4738
rect -8362 -100 -7296 1458
rect 32552 1424 32992 1952
rect 67046 1476 67496 1918
rect 13690 -202 14226 56
rect 48476 -266 48970 -26
rect -8406 -6996 -7286 -5478
rect 32570 -2002 33010 -1474
rect 68986 -1972 69404 -1496
rect 30 -4796 440 -4324
rect 34736 -4796 35036 -4302
rect 68986 -4784 69424 -4296
rect 30208 -5896 30568 -5580
rect 64870 -6024 65252 -5584
rect 82 -8234 432 -7728
rect 34740 -8240 35126 -7758
rect 66992 -8242 67518 -7724
rect -22 -11212 344 -10754
rect 34652 -11260 35046 -10764
rect -48 -14682 294 -14180
rect 34642 -14672 35026 -14192
rect 34608 -17502 35046 -16998
rect 13674 -18910 14250 -18696
rect 48494 -18870 48944 -18612
<< metal3 >>
rect 34608 8322 35192 8327
rect 34 8190 464 8195
rect 34 7678 44 8190
rect 454 7678 464 8190
rect 34 7673 464 7678
rect 34608 7624 34618 8322
rect 35182 7624 35192 8322
rect 68952 8282 69406 8287
rect 68952 7730 68962 8282
rect 69396 7730 69406 8282
rect 68952 7725 69406 7730
rect 34608 7619 35192 7624
rect 64872 5869 65238 5871
rect 64870 5866 65252 5869
rect 30208 5849 30564 5862
rect 30208 5844 30574 5849
rect 30208 5550 30222 5844
rect 30564 5550 30574 5844
rect 30208 5545 30574 5550
rect 64870 5550 64882 5866
rect 65228 5550 65252 5866
rect -3658 4731 374 4734
rect -3658 4726 454 4731
rect -3658 4240 28 4726
rect 444 4240 454 4726
rect -3658 4235 454 4240
rect -3658 4222 374 4235
rect -8372 1458 -7286 1463
rect -8372 -100 -8362 1458
rect -7296 -100 -7286 1458
rect -8372 -105 -7286 -100
rect -3650 -4316 -2690 4222
rect 13680 56 14236 61
rect 13680 -202 13690 56
rect 14226 -202 14236 56
rect 13680 -207 14236 -202
rect -3650 -4319 422 -4316
rect -3650 -4324 450 -4319
rect -3650 -4778 30 -4324
rect -8416 -5478 -7276 -5473
rect -8416 -6996 -8406 -5478
rect -7286 -5718 -7276 -5478
rect -3650 -5718 -2690 -4778
rect 20 -4796 30 -4778
rect 440 -4796 450 -4324
rect 20 -4801 450 -4796
rect 30208 -5575 30564 5545
rect 34714 4734 35132 4739
rect 34714 4721 34724 4734
rect 31731 4235 34724 4721
rect 31731 -4365 32061 4235
rect 34714 4230 34724 4235
rect 35122 4230 35132 4734
rect 34714 4225 35132 4230
rect 32542 1952 33002 1957
rect 32542 1424 32552 1952
rect 32992 1424 33002 1952
rect 32542 1419 33002 1424
rect 48466 -26 48980 -21
rect 48466 -266 48476 -26
rect 48970 -266 48980 -26
rect 48466 -271 48980 -266
rect 32560 -1474 33020 -1469
rect 32560 -2002 32570 -1474
rect 33010 -2002 33020 -1474
rect 32560 -2007 33020 -2002
rect 34726 -4302 35046 -4297
rect 34726 -4365 34736 -4302
rect 31731 -4773 34736 -4365
rect -7286 -6760 -2690 -5718
rect 30198 -5580 30578 -5575
rect 30198 -5896 30208 -5580
rect 30568 -5896 30578 -5580
rect 30198 -5901 30578 -5896
rect -7286 -6996 -7276 -6760
rect -8416 -7001 -7276 -6996
rect -3650 -14196 -2690 -6760
rect 72 -7728 442 -7723
rect 72 -8234 82 -7728
rect 432 -8234 442 -7728
rect 72 -8239 442 -8234
rect 30790 -8428 30800 -7702
rect 31198 -7836 31208 -7702
rect 31731 -7836 32061 -4773
rect 34726 -4796 34736 -4773
rect 35036 -4796 35046 -4302
rect 34726 -4801 35046 -4796
rect 64870 -5579 65252 5550
rect 68966 4738 69424 4743
rect 68966 4698 68976 4738
rect 66018 4322 68976 4698
rect 66018 -4380 66394 4322
rect 68966 4250 68976 4322
rect 69414 4250 69424 4738
rect 68966 4245 69424 4250
rect 67036 1918 67506 1923
rect 67036 1476 67046 1918
rect 67496 1476 67506 1918
rect 67036 1471 67506 1476
rect 68976 -1496 69414 -1491
rect 68976 -1972 68986 -1496
rect 69404 -1972 69414 -1496
rect 68976 -1977 69414 -1972
rect 68976 -4296 69434 -4291
rect 68976 -4380 68986 -4296
rect 66018 -4756 68986 -4380
rect 64860 -5584 65262 -5579
rect 64860 -6024 64870 -5584
rect 65252 -6024 65262 -5584
rect 64860 -6029 65262 -6024
rect 31198 -8270 32061 -7836
rect 34730 -7758 35136 -7753
rect 34730 -8240 34740 -7758
rect 35126 -8240 35136 -7758
rect 66018 -7824 66394 -4756
rect 68976 -4784 68986 -4756
rect 69424 -4784 69434 -4296
rect 68976 -4789 69434 -4784
rect 65498 -7832 66394 -7824
rect 34730 -8245 35136 -8240
rect 31198 -8428 31208 -8270
rect -32 -10754 354 -10749
rect -32 -11212 -22 -10754
rect 344 -11212 354 -10754
rect -32 -11217 354 -11212
rect -58 -14180 304 -14175
rect -58 -14196 -48 -14180
rect -3650 -14682 -48 -14196
rect 294 -14196 304 -14180
rect 294 -14682 330 -14196
rect 31731 -14211 32061 -8270
rect 65488 -8298 65498 -7832
rect 65830 -8298 66394 -7832
rect 66982 -7724 67528 -7719
rect 66982 -8242 66992 -7724
rect 67518 -8242 67528 -7724
rect 66982 -8247 67528 -8242
rect 34642 -10764 35056 -10759
rect 34642 -11260 34652 -10764
rect 35046 -11260 35056 -10764
rect 34642 -11265 35056 -11260
rect 34632 -14192 35036 -14187
rect 34632 -14211 34642 -14192
rect 31731 -14647 34642 -14211
rect 34632 -14672 34642 -14647
rect 35026 -14672 35036 -14192
rect 34632 -14677 35036 -14672
rect -3650 -14888 -2690 -14682
rect -58 -14687 304 -14682
rect 34598 -16998 35056 -16993
rect 34598 -17502 34608 -16998
rect 35046 -17502 35056 -16998
rect 34598 -17507 35056 -17502
rect 48484 -18612 48954 -18607
rect 13664 -18696 14260 -18691
rect 13664 -18910 13674 -18696
rect 14250 -18910 14260 -18696
rect 48484 -18870 48494 -18612
rect 48944 -18870 48954 -18612
rect 48484 -18875 48954 -18870
rect 13664 -18915 14260 -18910
<< via3 >>
rect 44 7678 454 8190
rect 34618 7624 35182 8322
rect 68962 7730 69396 8282
rect -8362 -100 -7296 1458
rect 13690 -202 14226 56
rect 32552 1424 32992 1952
rect 48476 -266 48970 -26
rect 32570 -2002 33010 -1474
rect 82 -8234 432 -7728
rect 30800 -8428 31198 -7702
rect 67046 1476 67496 1918
rect 68986 -1972 69404 -1496
rect 34740 -8240 35126 -7758
rect -22 -11212 344 -10754
rect 65498 -8298 65830 -7832
rect 66992 -8242 67518 -7724
rect 34652 -11260 35046 -10764
rect 34608 -17502 35046 -16998
rect 13674 -18910 14250 -18696
rect 48494 -18870 48944 -18612
<< metal4 >>
rect 34617 8322 35183 8323
rect 34617 8232 34618 8322
rect 43 8190 455 8191
rect 43 8168 44 8190
rect -1944 8139 44 8168
rect -1945 7706 44 8139
rect -8363 1458 -7295 1459
rect -8363 -100 -8362 1458
rect -7296 1170 -7295 1458
rect -1945 1170 -959 7706
rect 43 7678 44 7706
rect 454 8168 455 8190
rect 454 7706 461 8168
rect 30744 7770 34618 8232
rect 454 7678 455 7706
rect 43 7677 455 7678
rect 32562 1953 33002 1966
rect 32551 1952 33002 1953
rect 32551 1424 32552 1952
rect 32992 1424 33002 1952
rect 32551 1423 33002 1424
rect -7296 120 -959 1170
rect -7296 106 -6654 120
rect -7296 -100 -7295 106
rect -8363 -101 -7295 -100
rect -1945 -1494 -959 120
rect 13689 56 14227 57
rect 13689 -202 13690 56
rect 14226 -202 14227 56
rect 13689 -203 14227 -202
rect 32562 -1473 33002 1423
rect 32562 -1474 33011 -1473
rect -1945 -1974 -956 -1494
rect -1945 -7746 -959 -1974
rect 32562 -2002 32570 -1474
rect 33010 -2002 33011 -1474
rect 32562 -2003 33011 -2002
rect 30799 -7702 31199 -7701
rect 81 -7728 433 -7727
rect 81 -7746 82 -7728
rect -1945 -8234 82 -7746
rect 432 -8234 433 -7728
rect -1945 -8235 433 -8234
rect -1945 -8252 424 -8235
rect -1945 -10754 -959 -8252
rect 30799 -8428 30800 -7702
rect 31198 -8428 31199 -7702
rect 30799 -8429 31199 -8428
rect 32562 -10702 33002 -2003
rect -23 -10754 345 -10753
rect -1945 -11212 -22 -10754
rect 344 -11212 368 -10754
rect 30724 -11170 33002 -10702
rect -1945 -11244 368 -11212
rect -1945 -11349 -959 -11244
rect 32562 -17048 33002 -11170
rect 33501 -7779 33963 7770
rect 34617 7624 34618 7770
rect 35182 7624 35183 8322
rect 68961 8282 69397 8283
rect 68961 8230 68962 8282
rect 65430 7768 68962 8230
rect 34617 7623 35183 7624
rect 67039 1918 67501 2069
rect 67039 1476 67046 1918
rect 67496 1476 67501 1918
rect 48475 -266 48476 -260
rect 48970 -266 48971 -260
rect 48475 -267 48971 -266
rect 67039 -7723 67501 1476
rect 68099 -1481 68561 7768
rect 68961 7730 68962 7768
rect 69396 7730 69397 8282
rect 68961 7729 69397 7730
rect 99684 2343 100146 8234
rect 101138 2343 102002 3218
rect 99684 1881 102002 2343
rect 101138 1068 102002 1881
rect 68099 -1495 69367 -1481
rect 68099 -1496 69405 -1495
rect 68099 -1943 68986 -1496
rect 68985 -1972 68986 -1943
rect 69404 -1972 69405 -1496
rect 68985 -1973 69405 -1972
rect 66991 -7724 67519 -7723
rect 34739 -7758 35127 -7757
rect 34739 -7779 34740 -7758
rect 33501 -8240 34740 -7779
rect 35126 -8240 35127 -7758
rect 33501 -8241 35127 -8240
rect 65497 -7832 65831 -7831
rect 33501 -10785 33963 -8241
rect 65497 -8298 65498 -7832
rect 65830 -8298 65831 -7832
rect 66991 -8242 66992 -7724
rect 67518 -8242 67519 -7724
rect 101154 -7811 102018 -7008
rect 66991 -8243 67519 -8242
rect 65497 -8299 65831 -8298
rect 67039 -10696 67501 -8243
rect 99678 -8273 102018 -7811
rect 101154 -9158 102018 -8273
rect 34651 -10764 35047 -10763
rect 34651 -10785 34652 -10764
rect 33501 -11247 34652 -10785
rect 34651 -11260 34652 -11247
rect 35046 -11260 35047 -10764
rect 65334 -11158 67663 -10696
rect 34651 -11261 35047 -11260
rect 34607 -16998 35047 -16997
rect 34607 -17048 34608 -16998
rect 32562 -17488 34608 -17048
rect 34607 -17502 34608 -17488
rect 35046 -17502 35047 -16998
rect 34607 -17503 35047 -17502
rect 13673 -18696 13684 -18695
rect 48493 -18612 48945 -18611
rect 14224 -18696 14251 -18695
rect 13673 -18910 13674 -18696
rect 14250 -18910 14251 -18696
rect 48493 -18870 48494 -18612
rect 48944 -18870 48945 -18612
rect 48493 -18871 48945 -18870
rect 13673 -18911 14251 -18910
<< via4 >>
rect 13690 -202 14226 56
rect 48472 -26 48974 -16
rect 48472 -260 48476 -26
rect 48476 -260 48970 -26
rect 48970 -260 48974 -26
rect 13684 -18696 14224 -18550
rect 13684 -18888 14224 -18696
rect 48494 -18870 48944 -18612
<< metal5 >>
rect 13662 56 14254 100
rect 13662 -202 13690 56
rect 14226 -202 14254 56
rect 13662 -382 14254 -202
rect 48444 -16 49002 10
rect 48444 -260 48472 -16
rect 48974 -260 49002 -16
rect 48444 -362 49002 -260
rect 13674 -18526 14244 -382
rect 13660 -18550 14248 -18526
rect 13660 -18888 13684 -18550
rect 14224 -18888 14248 -18550
rect 48452 -18612 48996 -362
rect 48452 -18672 48494 -18612
rect 13660 -18912 14248 -18888
rect 48454 -18870 48494 -18672
rect 48944 -18672 48996 -18612
rect 48944 -18870 48994 -18672
rect 48454 -18904 48994 -18870
use analog_neuron_3input_re  analog_neuron_3input_re_0
timestamp 1627890010
transform 1 0 548 0 1 6266
box -548 -6266 30658 3151
use analog_neuron_3input_re  analog_neuron_3input_re_1
timestamp 1627890010
transform 1 0 550 0 -1 -6309
box -548 -6266 30658 3151
use analog_neuron_3input_re  analog_neuron_3input_re_2
timestamp 1627890010
transform 1 0 460 0 1 -12660
box -548 -6266 30658 3151
use analog_neuron_3input_re  analog_neuron_3input_re_3
timestamp 1627890010
transform 1 0 35234 0 1 6264
box -548 -6266 30658 3151
use analog_neuron_3input_re  analog_neuron_3input_re_4
timestamp 1627890010
transform 1 0 35236 0 -1 -6311
box -548 -6266 30658 3151
use analog_neuron_3input_re  analog_neuron_3input_re_5
timestamp 1627890010
transform 1 0 35146 0 1 -12662
box -548 -6266 30658 3151
use analog_neuron_3input_re  analog_neuron_3input_re_6
timestamp 1627890010
transform 1 0 69488 0 1 6268
box -548 -6266 30658 3151
use analog_neuron_3input_re  analog_neuron_3input_re_7
timestamp 1627890010
transform 1 0 69490 0 -1 -6307
box -548 -6266 30658 3151
<< labels >>
rlabel metal4 101282 -9094 101942 -7102 1 Out2
port 1 n
rlabel metal4 101208 1120 101868 3112 1 Out1
port 2 n
rlabel metal2 -8490 -382 -7204 1836 1 In1
port 3 n
rlabel metal2 -8528 -7322 -7242 -5104 1 In2
port 4 n
rlabel metal2 -8472 -13574 -7186 -11356 1 In3
port 5 n
rlabel metal2 1472 9288 99492 9404 1 VDD
port 6 n
rlabel metal2 2048 -18912 63536 -18810 1 GND
port 7 n
rlabel metal2 21232 -132 54090 64 1 GND
port 7 n
rlabel metal2 55578 -140 88294 60 1 GND
port 7 n
rlabel metal2 89822 -154 97866 90 1 GND
port 7 n
rlabel metal2 4408 -9582 36564 -9412 1 VDD
port 6 n
rlabel metal2 38920 -9594 99424 -9412 1 VDD
port 6 n
rlabel metal2 2040 -138 19166 102 1 GND
port 7 n
<< end >>
