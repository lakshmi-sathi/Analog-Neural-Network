magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< error_p >>
rect -29 -307 29 -301
rect -29 -341 -17 -307
rect -29 -347 29 -341
<< pwell >>
rect -175 409 175 443
rect -175 -409 -141 409
rect 141 -409 175 409
rect -175 -443 175 -409
<< nmos >>
rect -15 -269 15 331
<< ndiff >>
rect -73 286 -15 331
rect -73 252 -61 286
rect -27 252 -15 286
rect -73 218 -15 252
rect -73 184 -61 218
rect -27 184 -15 218
rect -73 150 -15 184
rect -73 116 -61 150
rect -27 116 -15 150
rect -73 82 -15 116
rect -73 48 -61 82
rect -27 48 -15 82
rect -73 14 -15 48
rect -73 -20 -61 14
rect -27 -20 -15 14
rect -73 -54 -15 -20
rect -73 -88 -61 -54
rect -27 -88 -15 -54
rect -73 -122 -15 -88
rect -73 -156 -61 -122
rect -27 -156 -15 -122
rect -73 -190 -15 -156
rect -73 -224 -61 -190
rect -27 -224 -15 -190
rect -73 -269 -15 -224
rect 15 286 73 331
rect 15 252 27 286
rect 61 252 73 286
rect 15 218 73 252
rect 15 184 27 218
rect 61 184 73 218
rect 15 150 73 184
rect 15 116 27 150
rect 61 116 73 150
rect 15 82 73 116
rect 15 48 27 82
rect 61 48 73 82
rect 15 14 73 48
rect 15 -20 27 14
rect 61 -20 73 14
rect 15 -54 73 -20
rect 15 -88 27 -54
rect 61 -88 73 -54
rect 15 -122 73 -88
rect 15 -156 27 -122
rect 61 -156 73 -122
rect 15 -190 73 -156
rect 15 -224 27 -190
rect 61 -224 73 -190
rect 15 -269 73 -224
<< ndiffc >>
rect -61 252 -27 286
rect -61 184 -27 218
rect -61 116 -27 150
rect -61 48 -27 82
rect -61 -20 -27 14
rect -61 -88 -27 -54
rect -61 -156 -27 -122
rect -61 -224 -27 -190
rect 27 252 61 286
rect 27 184 61 218
rect 27 116 61 150
rect 27 48 61 82
rect 27 -20 61 14
rect 27 -88 61 -54
rect 27 -156 61 -122
rect 27 -224 61 -190
<< psubdiff >>
rect -175 409 -51 443
rect -17 409 17 443
rect 51 409 175 443
rect -175 323 -141 409
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect 141 323 175 409
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect -175 -409 -141 -323
rect 141 -409 175 -323
rect -175 -443 -51 -409
rect -17 -443 17 -409
rect 51 -443 175 -409
<< psubdiffcont >>
rect -51 409 -17 443
rect 17 409 51 443
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect -175 -323 -141 -289
rect 141 -323 175 -289
rect -51 -443 -17 -409
rect 17 -443 51 -409
<< poly >>
rect -15 331 15 357
rect -15 -291 15 -269
rect -33 -307 33 -291
rect -33 -341 -17 -307
rect 17 -341 33 -307
rect -33 -357 33 -341
<< polycont >>
rect -17 -341 17 -307
<< locali >>
rect -175 409 -51 443
rect -17 409 17 443
rect 51 409 175 443
rect -175 323 -141 409
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect -61 300 -27 335
rect -61 228 -27 252
rect -61 156 -27 184
rect -61 84 -27 116
rect -61 14 -27 48
rect -61 -54 -27 -22
rect -61 -122 -27 -94
rect -61 -190 -27 -166
rect -61 -273 -27 -238
rect 27 300 61 335
rect 27 228 61 252
rect 27 156 61 184
rect 27 84 61 116
rect 27 14 61 48
rect 27 -54 61 -22
rect 27 -122 61 -94
rect 27 -190 61 -166
rect 27 -273 61 -238
rect 141 323 175 409
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect -175 -409 -141 -323
rect -33 -341 -17 -307
rect 17 -341 33 -307
rect 141 -409 175 -323
rect -175 -443 -51 -409
rect -17 -443 17 -409
rect 51 -443 175 -409
<< viali >>
rect -61 286 -27 300
rect -61 266 -27 286
rect -61 218 -27 228
rect -61 194 -27 218
rect -61 150 -27 156
rect -61 122 -27 150
rect -61 82 -27 84
rect -61 50 -27 82
rect -61 -20 -27 12
rect -61 -22 -27 -20
rect -61 -88 -27 -60
rect -61 -94 -27 -88
rect -61 -156 -27 -132
rect -61 -166 -27 -156
rect -61 -224 -27 -204
rect -61 -238 -27 -224
rect 27 286 61 300
rect 27 266 61 286
rect 27 218 61 228
rect 27 194 61 218
rect 27 150 61 156
rect 27 122 61 150
rect 27 82 61 84
rect 27 50 61 82
rect 27 -20 61 12
rect 27 -22 61 -20
rect 27 -88 61 -60
rect 27 -94 61 -88
rect 27 -156 61 -132
rect 27 -166 61 -156
rect 27 -224 61 -204
rect 27 -238 61 -224
rect -17 -341 17 -307
<< metal1 >>
rect -67 300 -21 331
rect -67 266 -61 300
rect -27 266 -21 300
rect -67 228 -21 266
rect -67 194 -61 228
rect -27 194 -21 228
rect -67 156 -21 194
rect -67 122 -61 156
rect -27 122 -21 156
rect -67 84 -21 122
rect -67 50 -61 84
rect -27 50 -21 84
rect -67 12 -21 50
rect -67 -22 -61 12
rect -27 -22 -21 12
rect -67 -60 -21 -22
rect -67 -94 -61 -60
rect -27 -94 -21 -60
rect -67 -132 -21 -94
rect -67 -166 -61 -132
rect -27 -166 -21 -132
rect -67 -204 -21 -166
rect -67 -238 -61 -204
rect -27 -238 -21 -204
rect -67 -269 -21 -238
rect 21 300 67 331
rect 21 266 27 300
rect 61 266 67 300
rect 21 228 67 266
rect 21 194 27 228
rect 61 194 67 228
rect 21 156 67 194
rect 21 122 27 156
rect 61 122 67 156
rect 21 84 67 122
rect 21 50 27 84
rect 61 50 67 84
rect 21 12 67 50
rect 21 -22 27 12
rect 61 -22 67 12
rect 21 -60 67 -22
rect 21 -94 27 -60
rect 61 -94 67 -60
rect 21 -132 67 -94
rect 21 -166 27 -132
rect 61 -166 67 -132
rect 21 -204 67 -166
rect 21 -238 27 -204
rect 61 -238 67 -204
rect 21 -269 67 -238
rect -29 -307 29 -301
rect -29 -341 -17 -307
rect 17 -341 29 -307
rect -29 -347 29 -341
<< properties >>
string FIXED_BBOX -158 -426 158 426
<< end >>
