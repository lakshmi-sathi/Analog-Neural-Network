magic
tech sky130A
magscale 1 2
timestamp 1626793425
<< error_p >>
rect -1814 641 -1756 647
rect -1394 641 -1336 647
rect -974 641 -916 647
rect -554 641 -496 647
rect -134 641 -76 647
rect 286 641 344 647
rect 706 641 764 647
rect 1126 641 1184 647
rect 1546 641 1604 647
rect -1814 607 -1802 641
rect -1394 607 -1382 641
rect -974 607 -962 641
rect -554 607 -542 641
rect -134 607 -122 641
rect 286 607 298 641
rect 706 607 718 641
rect 1126 607 1138 641
rect 1546 607 1558 641
rect -1814 601 -1756 607
rect -1394 601 -1336 607
rect -974 601 -916 607
rect -554 601 -496 607
rect -134 601 -76 607
rect 286 601 344 607
rect 706 601 764 607
rect 1126 601 1184 607
rect 1546 601 1604 607
rect -1604 71 -1546 77
rect -1184 71 -1126 77
rect -764 71 -706 77
rect -344 71 -286 77
rect 76 71 134 77
rect 496 71 554 77
rect 916 71 974 77
rect 1336 71 1394 77
rect 1756 71 1814 77
rect -1604 37 -1592 71
rect -1184 37 -1172 71
rect -764 37 -752 71
rect -344 37 -332 71
rect 76 37 88 71
rect 496 37 508 71
rect 916 37 928 71
rect 1336 37 1348 71
rect 1756 37 1768 71
rect -1604 31 -1546 37
rect -1184 31 -1126 37
rect -764 31 -706 37
rect -344 31 -286 37
rect 76 31 134 37
rect 496 31 554 37
rect 916 31 974 37
rect 1336 31 1394 37
rect 1756 31 1814 37
rect -1604 -37 -1546 -31
rect -1184 -37 -1126 -31
rect -764 -37 -706 -31
rect -344 -37 -286 -31
rect 76 -37 134 -31
rect 496 -37 554 -31
rect 916 -37 974 -31
rect 1336 -37 1394 -31
rect 1756 -37 1814 -31
rect -1604 -71 -1592 -37
rect -1184 -71 -1172 -37
rect -764 -71 -752 -37
rect -344 -71 -332 -37
rect 76 -71 88 -37
rect 496 -71 508 -37
rect 916 -71 928 -37
rect 1336 -71 1348 -37
rect 1756 -71 1768 -37
rect -1604 -77 -1546 -71
rect -1184 -77 -1126 -71
rect -764 -77 -706 -71
rect -344 -77 -286 -71
rect 76 -77 134 -71
rect 496 -77 554 -71
rect 916 -77 974 -71
rect 1336 -77 1394 -71
rect 1756 -77 1814 -71
rect -1814 -607 -1756 -601
rect -1394 -607 -1336 -601
rect -974 -607 -916 -601
rect -554 -607 -496 -601
rect -134 -607 -76 -601
rect 286 -607 344 -601
rect 706 -607 764 -601
rect 1126 -607 1184 -601
rect 1546 -607 1604 -601
rect -1814 -641 -1802 -607
rect -1394 -641 -1382 -607
rect -974 -641 -962 -607
rect -554 -641 -542 -607
rect -134 -641 -122 -607
rect 286 -641 298 -607
rect 706 -641 718 -607
rect 1126 -641 1138 -607
rect 1546 -641 1558 -607
rect -1814 -647 -1756 -641
rect -1394 -647 -1336 -641
rect -974 -647 -916 -641
rect -554 -647 -496 -641
rect -134 -647 -76 -641
rect 286 -647 344 -641
rect 706 -647 764 -641
rect 1126 -647 1184 -641
rect 1546 -647 1604 -641
<< nwell >>
rect -2000 -779 2000 779
<< pmos >>
rect -1800 118 -1770 560
rect -1590 118 -1560 560
rect -1380 118 -1350 560
rect -1170 118 -1140 560
rect -960 118 -930 560
rect -750 118 -720 560
rect -540 118 -510 560
rect -330 118 -300 560
rect -120 118 -90 560
rect 90 118 120 560
rect 300 118 330 560
rect 510 118 540 560
rect 720 118 750 560
rect 930 118 960 560
rect 1140 118 1170 560
rect 1350 118 1380 560
rect 1560 118 1590 560
rect 1770 118 1800 560
rect -1800 -560 -1770 -118
rect -1590 -560 -1560 -118
rect -1380 -560 -1350 -118
rect -1170 -560 -1140 -118
rect -960 -560 -930 -118
rect -750 -560 -720 -118
rect -540 -560 -510 -118
rect -330 -560 -300 -118
rect -120 -560 -90 -118
rect 90 -560 120 -118
rect 300 -560 330 -118
rect 510 -560 540 -118
rect 720 -560 750 -118
rect 930 -560 960 -118
rect 1140 -560 1170 -118
rect 1350 -560 1380 -118
rect 1560 -560 1590 -118
rect 1770 -560 1800 -118
<< pdiff >>
rect -1862 548 -1800 560
rect -1862 130 -1850 548
rect -1816 130 -1800 548
rect -1862 118 -1800 130
rect -1770 548 -1708 560
rect -1770 130 -1754 548
rect -1720 130 -1708 548
rect -1770 118 -1708 130
rect -1652 548 -1590 560
rect -1652 130 -1640 548
rect -1606 130 -1590 548
rect -1652 118 -1590 130
rect -1560 548 -1498 560
rect -1560 130 -1544 548
rect -1510 130 -1498 548
rect -1560 118 -1498 130
rect -1442 548 -1380 560
rect -1442 130 -1430 548
rect -1396 130 -1380 548
rect -1442 118 -1380 130
rect -1350 548 -1288 560
rect -1350 130 -1334 548
rect -1300 130 -1288 548
rect -1350 118 -1288 130
rect -1232 548 -1170 560
rect -1232 130 -1220 548
rect -1186 130 -1170 548
rect -1232 118 -1170 130
rect -1140 548 -1078 560
rect -1140 130 -1124 548
rect -1090 130 -1078 548
rect -1140 118 -1078 130
rect -1022 548 -960 560
rect -1022 130 -1010 548
rect -976 130 -960 548
rect -1022 118 -960 130
rect -930 548 -868 560
rect -930 130 -914 548
rect -880 130 -868 548
rect -930 118 -868 130
rect -812 548 -750 560
rect -812 130 -800 548
rect -766 130 -750 548
rect -812 118 -750 130
rect -720 548 -658 560
rect -720 130 -704 548
rect -670 130 -658 548
rect -720 118 -658 130
rect -602 548 -540 560
rect -602 130 -590 548
rect -556 130 -540 548
rect -602 118 -540 130
rect -510 548 -448 560
rect -510 130 -494 548
rect -460 130 -448 548
rect -510 118 -448 130
rect -392 548 -330 560
rect -392 130 -380 548
rect -346 130 -330 548
rect -392 118 -330 130
rect -300 548 -238 560
rect -300 130 -284 548
rect -250 130 -238 548
rect -300 118 -238 130
rect -182 548 -120 560
rect -182 130 -170 548
rect -136 130 -120 548
rect -182 118 -120 130
rect -90 548 -28 560
rect -90 130 -74 548
rect -40 130 -28 548
rect -90 118 -28 130
rect 28 548 90 560
rect 28 130 40 548
rect 74 130 90 548
rect 28 118 90 130
rect 120 548 182 560
rect 120 130 136 548
rect 170 130 182 548
rect 120 118 182 130
rect 238 548 300 560
rect 238 130 250 548
rect 284 130 300 548
rect 238 118 300 130
rect 330 548 392 560
rect 330 130 346 548
rect 380 130 392 548
rect 330 118 392 130
rect 448 548 510 560
rect 448 130 460 548
rect 494 130 510 548
rect 448 118 510 130
rect 540 548 602 560
rect 540 130 556 548
rect 590 130 602 548
rect 540 118 602 130
rect 658 548 720 560
rect 658 130 670 548
rect 704 130 720 548
rect 658 118 720 130
rect 750 548 812 560
rect 750 130 766 548
rect 800 130 812 548
rect 750 118 812 130
rect 868 548 930 560
rect 868 130 880 548
rect 914 130 930 548
rect 868 118 930 130
rect 960 548 1022 560
rect 960 130 976 548
rect 1010 130 1022 548
rect 960 118 1022 130
rect 1078 548 1140 560
rect 1078 130 1090 548
rect 1124 130 1140 548
rect 1078 118 1140 130
rect 1170 548 1232 560
rect 1170 130 1186 548
rect 1220 130 1232 548
rect 1170 118 1232 130
rect 1288 548 1350 560
rect 1288 130 1300 548
rect 1334 130 1350 548
rect 1288 118 1350 130
rect 1380 548 1442 560
rect 1380 130 1396 548
rect 1430 130 1442 548
rect 1380 118 1442 130
rect 1498 548 1560 560
rect 1498 130 1510 548
rect 1544 130 1560 548
rect 1498 118 1560 130
rect 1590 548 1652 560
rect 1590 130 1606 548
rect 1640 130 1652 548
rect 1590 118 1652 130
rect 1708 548 1770 560
rect 1708 130 1720 548
rect 1754 130 1770 548
rect 1708 118 1770 130
rect 1800 548 1862 560
rect 1800 130 1816 548
rect 1850 130 1862 548
rect 1800 118 1862 130
rect -1862 -130 -1800 -118
rect -1862 -548 -1850 -130
rect -1816 -548 -1800 -130
rect -1862 -560 -1800 -548
rect -1770 -130 -1708 -118
rect -1770 -548 -1754 -130
rect -1720 -548 -1708 -130
rect -1770 -560 -1708 -548
rect -1652 -130 -1590 -118
rect -1652 -548 -1640 -130
rect -1606 -548 -1590 -130
rect -1652 -560 -1590 -548
rect -1560 -130 -1498 -118
rect -1560 -548 -1544 -130
rect -1510 -548 -1498 -130
rect -1560 -560 -1498 -548
rect -1442 -130 -1380 -118
rect -1442 -548 -1430 -130
rect -1396 -548 -1380 -130
rect -1442 -560 -1380 -548
rect -1350 -130 -1288 -118
rect -1350 -548 -1334 -130
rect -1300 -548 -1288 -130
rect -1350 -560 -1288 -548
rect -1232 -130 -1170 -118
rect -1232 -548 -1220 -130
rect -1186 -548 -1170 -130
rect -1232 -560 -1170 -548
rect -1140 -130 -1078 -118
rect -1140 -548 -1124 -130
rect -1090 -548 -1078 -130
rect -1140 -560 -1078 -548
rect -1022 -130 -960 -118
rect -1022 -548 -1010 -130
rect -976 -548 -960 -130
rect -1022 -560 -960 -548
rect -930 -130 -868 -118
rect -930 -548 -914 -130
rect -880 -548 -868 -130
rect -930 -560 -868 -548
rect -812 -130 -750 -118
rect -812 -548 -800 -130
rect -766 -548 -750 -130
rect -812 -560 -750 -548
rect -720 -130 -658 -118
rect -720 -548 -704 -130
rect -670 -548 -658 -130
rect -720 -560 -658 -548
rect -602 -130 -540 -118
rect -602 -548 -590 -130
rect -556 -548 -540 -130
rect -602 -560 -540 -548
rect -510 -130 -448 -118
rect -510 -548 -494 -130
rect -460 -548 -448 -130
rect -510 -560 -448 -548
rect -392 -130 -330 -118
rect -392 -548 -380 -130
rect -346 -548 -330 -130
rect -392 -560 -330 -548
rect -300 -130 -238 -118
rect -300 -548 -284 -130
rect -250 -548 -238 -130
rect -300 -560 -238 -548
rect -182 -130 -120 -118
rect -182 -548 -170 -130
rect -136 -548 -120 -130
rect -182 -560 -120 -548
rect -90 -130 -28 -118
rect -90 -548 -74 -130
rect -40 -548 -28 -130
rect -90 -560 -28 -548
rect 28 -130 90 -118
rect 28 -548 40 -130
rect 74 -548 90 -130
rect 28 -560 90 -548
rect 120 -130 182 -118
rect 120 -548 136 -130
rect 170 -548 182 -130
rect 120 -560 182 -548
rect 238 -130 300 -118
rect 238 -548 250 -130
rect 284 -548 300 -130
rect 238 -560 300 -548
rect 330 -130 392 -118
rect 330 -548 346 -130
rect 380 -548 392 -130
rect 330 -560 392 -548
rect 448 -130 510 -118
rect 448 -548 460 -130
rect 494 -548 510 -130
rect 448 -560 510 -548
rect 540 -130 602 -118
rect 540 -548 556 -130
rect 590 -548 602 -130
rect 540 -560 602 -548
rect 658 -130 720 -118
rect 658 -548 670 -130
rect 704 -548 720 -130
rect 658 -560 720 -548
rect 750 -130 812 -118
rect 750 -548 766 -130
rect 800 -548 812 -130
rect 750 -560 812 -548
rect 868 -130 930 -118
rect 868 -548 880 -130
rect 914 -548 930 -130
rect 868 -560 930 -548
rect 960 -130 1022 -118
rect 960 -548 976 -130
rect 1010 -548 1022 -130
rect 960 -560 1022 -548
rect 1078 -130 1140 -118
rect 1078 -548 1090 -130
rect 1124 -548 1140 -130
rect 1078 -560 1140 -548
rect 1170 -130 1232 -118
rect 1170 -548 1186 -130
rect 1220 -548 1232 -130
rect 1170 -560 1232 -548
rect 1288 -130 1350 -118
rect 1288 -548 1300 -130
rect 1334 -548 1350 -130
rect 1288 -560 1350 -548
rect 1380 -130 1442 -118
rect 1380 -548 1396 -130
rect 1430 -548 1442 -130
rect 1380 -560 1442 -548
rect 1498 -130 1560 -118
rect 1498 -548 1510 -130
rect 1544 -548 1560 -130
rect 1498 -560 1560 -548
rect 1590 -130 1652 -118
rect 1590 -548 1606 -130
rect 1640 -548 1652 -130
rect 1590 -560 1652 -548
rect 1708 -130 1770 -118
rect 1708 -548 1720 -130
rect 1754 -548 1770 -130
rect 1708 -560 1770 -548
rect 1800 -130 1862 -118
rect 1800 -548 1816 -130
rect 1850 -548 1862 -130
rect 1800 -560 1862 -548
<< pdiffc >>
rect -1850 130 -1816 548
rect -1754 130 -1720 548
rect -1640 130 -1606 548
rect -1544 130 -1510 548
rect -1430 130 -1396 548
rect -1334 130 -1300 548
rect -1220 130 -1186 548
rect -1124 130 -1090 548
rect -1010 130 -976 548
rect -914 130 -880 548
rect -800 130 -766 548
rect -704 130 -670 548
rect -590 130 -556 548
rect -494 130 -460 548
rect -380 130 -346 548
rect -284 130 -250 548
rect -170 130 -136 548
rect -74 130 -40 548
rect 40 130 74 548
rect 136 130 170 548
rect 250 130 284 548
rect 346 130 380 548
rect 460 130 494 548
rect 556 130 590 548
rect 670 130 704 548
rect 766 130 800 548
rect 880 130 914 548
rect 976 130 1010 548
rect 1090 130 1124 548
rect 1186 130 1220 548
rect 1300 130 1334 548
rect 1396 130 1430 548
rect 1510 130 1544 548
rect 1606 130 1640 548
rect 1720 130 1754 548
rect 1816 130 1850 548
rect -1850 -548 -1816 -130
rect -1754 -548 -1720 -130
rect -1640 -548 -1606 -130
rect -1544 -548 -1510 -130
rect -1430 -548 -1396 -130
rect -1334 -548 -1300 -130
rect -1220 -548 -1186 -130
rect -1124 -548 -1090 -130
rect -1010 -548 -976 -130
rect -914 -548 -880 -130
rect -800 -548 -766 -130
rect -704 -548 -670 -130
rect -590 -548 -556 -130
rect -494 -548 -460 -130
rect -380 -548 -346 -130
rect -284 -548 -250 -130
rect -170 -548 -136 -130
rect -74 -548 -40 -130
rect 40 -548 74 -130
rect 136 -548 170 -130
rect 250 -548 284 -130
rect 346 -548 380 -130
rect 460 -548 494 -130
rect 556 -548 590 -130
rect 670 -548 704 -130
rect 766 -548 800 -130
rect 880 -548 914 -130
rect 976 -548 1010 -130
rect 1090 -548 1124 -130
rect 1186 -548 1220 -130
rect 1300 -548 1334 -130
rect 1396 -548 1430 -130
rect 1510 -548 1544 -130
rect 1606 -548 1640 -130
rect 1720 -548 1754 -130
rect 1816 -548 1850 -130
<< nsubdiff >>
rect -1964 709 -1868 743
rect 1868 709 1964 743
rect -1964 647 -1930 709
rect 1930 647 1964 709
rect -1964 -709 -1930 -647
rect 1930 -709 1964 -647
rect -1964 -743 -1868 -709
rect 1868 -743 1964 -709
<< nsubdiffcont >>
rect -1868 709 1868 743
rect -1964 -647 -1930 647
rect 1930 -647 1964 647
rect -1868 -743 1868 -709
<< poly >>
rect -1818 641 -1752 657
rect -1818 607 -1802 641
rect -1768 607 -1752 641
rect -1818 591 -1752 607
rect -1398 641 -1332 657
rect -1398 607 -1382 641
rect -1348 607 -1332 641
rect -1398 591 -1332 607
rect -978 641 -912 657
rect -978 607 -962 641
rect -928 607 -912 641
rect -978 591 -912 607
rect -558 641 -492 657
rect -558 607 -542 641
rect -508 607 -492 641
rect -558 591 -492 607
rect -138 641 -72 657
rect -138 607 -122 641
rect -88 607 -72 641
rect -138 591 -72 607
rect 282 641 348 657
rect 282 607 298 641
rect 332 607 348 641
rect 282 591 348 607
rect 702 641 768 657
rect 702 607 718 641
rect 752 607 768 641
rect 702 591 768 607
rect 1122 641 1188 657
rect 1122 607 1138 641
rect 1172 607 1188 641
rect 1122 591 1188 607
rect 1542 641 1608 657
rect 1542 607 1558 641
rect 1592 607 1608 641
rect 1542 591 1608 607
rect -1800 560 -1770 591
rect -1590 560 -1560 586
rect -1380 560 -1350 591
rect -1170 560 -1140 586
rect -960 560 -930 591
rect -750 560 -720 586
rect -540 560 -510 591
rect -330 560 -300 586
rect -120 560 -90 591
rect 90 560 120 586
rect 300 560 330 591
rect 510 560 540 586
rect 720 560 750 591
rect 930 560 960 586
rect 1140 560 1170 591
rect 1350 560 1380 586
rect 1560 560 1590 591
rect 1770 560 1800 586
rect -1800 92 -1770 118
rect -1590 87 -1560 118
rect -1380 92 -1350 118
rect -1170 87 -1140 118
rect -960 92 -930 118
rect -750 87 -720 118
rect -540 92 -510 118
rect -330 87 -300 118
rect -120 92 -90 118
rect 90 87 120 118
rect 300 92 330 118
rect 510 87 540 118
rect 720 92 750 118
rect 930 87 960 118
rect 1140 92 1170 118
rect 1350 87 1380 118
rect 1560 92 1590 118
rect 1770 87 1800 118
rect -1608 71 -1542 87
rect -1608 37 -1592 71
rect -1558 37 -1542 71
rect -1608 21 -1542 37
rect -1188 71 -1122 87
rect -1188 37 -1172 71
rect -1138 37 -1122 71
rect -1188 21 -1122 37
rect -768 71 -702 87
rect -768 37 -752 71
rect -718 37 -702 71
rect -768 21 -702 37
rect -348 71 -282 87
rect -348 37 -332 71
rect -298 37 -282 71
rect -348 21 -282 37
rect 72 71 138 87
rect 72 37 88 71
rect 122 37 138 71
rect 72 21 138 37
rect 492 71 558 87
rect 492 37 508 71
rect 542 37 558 71
rect 492 21 558 37
rect 912 71 978 87
rect 912 37 928 71
rect 962 37 978 71
rect 912 21 978 37
rect 1332 71 1398 87
rect 1332 37 1348 71
rect 1382 37 1398 71
rect 1332 21 1398 37
rect 1752 71 1818 87
rect 1752 37 1768 71
rect 1802 37 1818 71
rect 1752 21 1818 37
rect -1608 -37 -1542 -21
rect -1608 -71 -1592 -37
rect -1558 -71 -1542 -37
rect -1608 -87 -1542 -71
rect -1188 -37 -1122 -21
rect -1188 -71 -1172 -37
rect -1138 -71 -1122 -37
rect -1188 -87 -1122 -71
rect -768 -37 -702 -21
rect -768 -71 -752 -37
rect -718 -71 -702 -37
rect -768 -87 -702 -71
rect -348 -37 -282 -21
rect -348 -71 -332 -37
rect -298 -71 -282 -37
rect -348 -87 -282 -71
rect 72 -37 138 -21
rect 72 -71 88 -37
rect 122 -71 138 -37
rect 72 -87 138 -71
rect 492 -37 558 -21
rect 492 -71 508 -37
rect 542 -71 558 -37
rect 492 -87 558 -71
rect 912 -37 978 -21
rect 912 -71 928 -37
rect 962 -71 978 -37
rect 912 -87 978 -71
rect 1332 -37 1398 -21
rect 1332 -71 1348 -37
rect 1382 -71 1398 -37
rect 1332 -87 1398 -71
rect 1752 -37 1818 -21
rect 1752 -71 1768 -37
rect 1802 -71 1818 -37
rect 1752 -87 1818 -71
rect -1800 -118 -1770 -92
rect -1590 -118 -1560 -87
rect -1380 -118 -1350 -92
rect -1170 -118 -1140 -87
rect -960 -118 -930 -92
rect -750 -118 -720 -87
rect -540 -118 -510 -92
rect -330 -118 -300 -87
rect -120 -118 -90 -92
rect 90 -118 120 -87
rect 300 -118 330 -92
rect 510 -118 540 -87
rect 720 -118 750 -92
rect 930 -118 960 -87
rect 1140 -118 1170 -92
rect 1350 -118 1380 -87
rect 1560 -118 1590 -92
rect 1770 -118 1800 -87
rect -1800 -591 -1770 -560
rect -1590 -586 -1560 -560
rect -1380 -591 -1350 -560
rect -1170 -586 -1140 -560
rect -960 -591 -930 -560
rect -750 -586 -720 -560
rect -540 -591 -510 -560
rect -330 -586 -300 -560
rect -120 -591 -90 -560
rect 90 -586 120 -560
rect 300 -591 330 -560
rect 510 -586 540 -560
rect 720 -591 750 -560
rect 930 -586 960 -560
rect 1140 -591 1170 -560
rect 1350 -586 1380 -560
rect 1560 -591 1590 -560
rect 1770 -586 1800 -560
rect -1818 -607 -1752 -591
rect -1818 -641 -1802 -607
rect -1768 -641 -1752 -607
rect -1818 -657 -1752 -641
rect -1398 -607 -1332 -591
rect -1398 -641 -1382 -607
rect -1348 -641 -1332 -607
rect -1398 -657 -1332 -641
rect -978 -607 -912 -591
rect -978 -641 -962 -607
rect -928 -641 -912 -607
rect -978 -657 -912 -641
rect -558 -607 -492 -591
rect -558 -641 -542 -607
rect -508 -641 -492 -607
rect -558 -657 -492 -641
rect -138 -607 -72 -591
rect -138 -641 -122 -607
rect -88 -641 -72 -607
rect -138 -657 -72 -641
rect 282 -607 348 -591
rect 282 -641 298 -607
rect 332 -641 348 -607
rect 282 -657 348 -641
rect 702 -607 768 -591
rect 702 -641 718 -607
rect 752 -641 768 -607
rect 702 -657 768 -641
rect 1122 -607 1188 -591
rect 1122 -641 1138 -607
rect 1172 -641 1188 -607
rect 1122 -657 1188 -641
rect 1542 -607 1608 -591
rect 1542 -641 1558 -607
rect 1592 -641 1608 -607
rect 1542 -657 1608 -641
<< polycont >>
rect -1802 607 -1768 641
rect -1382 607 -1348 641
rect -962 607 -928 641
rect -542 607 -508 641
rect -122 607 -88 641
rect 298 607 332 641
rect 718 607 752 641
rect 1138 607 1172 641
rect 1558 607 1592 641
rect -1592 37 -1558 71
rect -1172 37 -1138 71
rect -752 37 -718 71
rect -332 37 -298 71
rect 88 37 122 71
rect 508 37 542 71
rect 928 37 962 71
rect 1348 37 1382 71
rect 1768 37 1802 71
rect -1592 -71 -1558 -37
rect -1172 -71 -1138 -37
rect -752 -71 -718 -37
rect -332 -71 -298 -37
rect 88 -71 122 -37
rect 508 -71 542 -37
rect 928 -71 962 -37
rect 1348 -71 1382 -37
rect 1768 -71 1802 -37
rect -1802 -641 -1768 -607
rect -1382 -641 -1348 -607
rect -962 -641 -928 -607
rect -542 -641 -508 -607
rect -122 -641 -88 -607
rect 298 -641 332 -607
rect 718 -641 752 -607
rect 1138 -641 1172 -607
rect 1558 -641 1592 -607
<< locali >>
rect -1964 709 -1868 743
rect 1868 709 1964 743
rect -1964 647 -1930 709
rect 1930 647 1964 709
rect -1818 607 -1802 641
rect -1768 607 -1752 641
rect -1398 607 -1382 641
rect -1348 607 -1332 641
rect -978 607 -962 641
rect -928 607 -912 641
rect -558 607 -542 641
rect -508 607 -492 641
rect -138 607 -122 641
rect -88 607 -72 641
rect 282 607 298 641
rect 332 607 348 641
rect 702 607 718 641
rect 752 607 768 641
rect 1122 607 1138 641
rect 1172 607 1188 641
rect 1542 607 1558 641
rect 1592 607 1608 641
rect -1850 548 -1816 564
rect -1850 114 -1816 130
rect -1754 548 -1720 564
rect -1754 114 -1720 130
rect -1640 548 -1606 564
rect -1640 114 -1606 130
rect -1544 548 -1510 564
rect -1544 114 -1510 130
rect -1430 548 -1396 564
rect -1430 114 -1396 130
rect -1334 548 -1300 564
rect -1334 114 -1300 130
rect -1220 548 -1186 564
rect -1220 114 -1186 130
rect -1124 548 -1090 564
rect -1124 114 -1090 130
rect -1010 548 -976 564
rect -1010 114 -976 130
rect -914 548 -880 564
rect -914 114 -880 130
rect -800 548 -766 564
rect -800 114 -766 130
rect -704 548 -670 564
rect -704 114 -670 130
rect -590 548 -556 564
rect -590 114 -556 130
rect -494 548 -460 564
rect -494 114 -460 130
rect -380 548 -346 564
rect -380 114 -346 130
rect -284 548 -250 564
rect -284 114 -250 130
rect -170 548 -136 564
rect -170 114 -136 130
rect -74 548 -40 564
rect -74 114 -40 130
rect 40 548 74 564
rect 40 114 74 130
rect 136 548 170 564
rect 136 114 170 130
rect 250 548 284 564
rect 250 114 284 130
rect 346 548 380 564
rect 346 114 380 130
rect 460 548 494 564
rect 460 114 494 130
rect 556 548 590 564
rect 556 114 590 130
rect 670 548 704 564
rect 670 114 704 130
rect 766 548 800 564
rect 766 114 800 130
rect 880 548 914 564
rect 880 114 914 130
rect 976 548 1010 564
rect 976 114 1010 130
rect 1090 548 1124 564
rect 1090 114 1124 130
rect 1186 548 1220 564
rect 1186 114 1220 130
rect 1300 548 1334 564
rect 1300 114 1334 130
rect 1396 548 1430 564
rect 1396 114 1430 130
rect 1510 548 1544 564
rect 1510 114 1544 130
rect 1606 548 1640 564
rect 1606 114 1640 130
rect 1720 548 1754 564
rect 1720 114 1754 130
rect 1816 548 1850 564
rect 1816 114 1850 130
rect -1608 37 -1592 71
rect -1558 37 -1542 71
rect -1188 37 -1172 71
rect -1138 37 -1122 71
rect -768 37 -752 71
rect -718 37 -702 71
rect -348 37 -332 71
rect -298 37 -282 71
rect 72 37 88 71
rect 122 37 138 71
rect 492 37 508 71
rect 542 37 558 71
rect 912 37 928 71
rect 962 37 978 71
rect 1332 37 1348 71
rect 1382 37 1398 71
rect 1752 37 1768 71
rect 1802 37 1818 71
rect -1608 -71 -1592 -37
rect -1558 -71 -1542 -37
rect -1188 -71 -1172 -37
rect -1138 -71 -1122 -37
rect -768 -71 -752 -37
rect -718 -71 -702 -37
rect -348 -71 -332 -37
rect -298 -71 -282 -37
rect 72 -71 88 -37
rect 122 -71 138 -37
rect 492 -71 508 -37
rect 542 -71 558 -37
rect 912 -71 928 -37
rect 962 -71 978 -37
rect 1332 -71 1348 -37
rect 1382 -71 1398 -37
rect 1752 -71 1768 -37
rect 1802 -71 1818 -37
rect -1850 -130 -1816 -114
rect -1850 -564 -1816 -548
rect -1754 -130 -1720 -114
rect -1754 -564 -1720 -548
rect -1640 -130 -1606 -114
rect -1640 -564 -1606 -548
rect -1544 -130 -1510 -114
rect -1544 -564 -1510 -548
rect -1430 -130 -1396 -114
rect -1430 -564 -1396 -548
rect -1334 -130 -1300 -114
rect -1334 -564 -1300 -548
rect -1220 -130 -1186 -114
rect -1220 -564 -1186 -548
rect -1124 -130 -1090 -114
rect -1124 -564 -1090 -548
rect -1010 -130 -976 -114
rect -1010 -564 -976 -548
rect -914 -130 -880 -114
rect -914 -564 -880 -548
rect -800 -130 -766 -114
rect -800 -564 -766 -548
rect -704 -130 -670 -114
rect -704 -564 -670 -548
rect -590 -130 -556 -114
rect -590 -564 -556 -548
rect -494 -130 -460 -114
rect -494 -564 -460 -548
rect -380 -130 -346 -114
rect -380 -564 -346 -548
rect -284 -130 -250 -114
rect -284 -564 -250 -548
rect -170 -130 -136 -114
rect -170 -564 -136 -548
rect -74 -130 -40 -114
rect -74 -564 -40 -548
rect 40 -130 74 -114
rect 40 -564 74 -548
rect 136 -130 170 -114
rect 136 -564 170 -548
rect 250 -130 284 -114
rect 250 -564 284 -548
rect 346 -130 380 -114
rect 346 -564 380 -548
rect 460 -130 494 -114
rect 460 -564 494 -548
rect 556 -130 590 -114
rect 556 -564 590 -548
rect 670 -130 704 -114
rect 670 -564 704 -548
rect 766 -130 800 -114
rect 766 -564 800 -548
rect 880 -130 914 -114
rect 880 -564 914 -548
rect 976 -130 1010 -114
rect 976 -564 1010 -548
rect 1090 -130 1124 -114
rect 1090 -564 1124 -548
rect 1186 -130 1220 -114
rect 1186 -564 1220 -548
rect 1300 -130 1334 -114
rect 1300 -564 1334 -548
rect 1396 -130 1430 -114
rect 1396 -564 1430 -548
rect 1510 -130 1544 -114
rect 1510 -564 1544 -548
rect 1606 -130 1640 -114
rect 1606 -564 1640 -548
rect 1720 -130 1754 -114
rect 1720 -564 1754 -548
rect 1816 -130 1850 -114
rect 1816 -564 1850 -548
rect -1818 -641 -1802 -607
rect -1768 -641 -1752 -607
rect -1398 -641 -1382 -607
rect -1348 -641 -1332 -607
rect -978 -641 -962 -607
rect -928 -641 -912 -607
rect -558 -641 -542 -607
rect -508 -641 -492 -607
rect -138 -641 -122 -607
rect -88 -641 -72 -607
rect 282 -641 298 -607
rect 332 -641 348 -607
rect 702 -641 718 -607
rect 752 -641 768 -607
rect 1122 -641 1138 -607
rect 1172 -641 1188 -607
rect 1542 -641 1558 -607
rect 1592 -641 1608 -607
rect -1964 -709 -1930 -647
rect 1930 -709 1964 -647
rect -1964 -743 -1868 -709
rect 1868 -743 1964 -709
<< viali >>
rect -1802 607 -1768 641
rect -1382 607 -1348 641
rect -962 607 -928 641
rect -542 607 -508 641
rect -122 607 -88 641
rect 298 607 332 641
rect 718 607 752 641
rect 1138 607 1172 641
rect 1558 607 1592 641
rect -1850 130 -1816 548
rect -1754 130 -1720 548
rect -1640 130 -1606 548
rect -1544 130 -1510 548
rect -1430 130 -1396 548
rect -1334 130 -1300 548
rect -1220 130 -1186 548
rect -1124 130 -1090 548
rect -1010 130 -976 548
rect -914 130 -880 548
rect -800 130 -766 548
rect -704 130 -670 548
rect -590 130 -556 548
rect -494 130 -460 548
rect -380 130 -346 548
rect -284 130 -250 548
rect -170 130 -136 548
rect -74 130 -40 548
rect 40 130 74 548
rect 136 130 170 548
rect 250 130 284 548
rect 346 130 380 548
rect 460 130 494 548
rect 556 130 590 548
rect 670 130 704 548
rect 766 130 800 548
rect 880 130 914 548
rect 976 130 1010 548
rect 1090 130 1124 548
rect 1186 130 1220 548
rect 1300 130 1334 548
rect 1396 130 1430 548
rect 1510 130 1544 548
rect 1606 130 1640 548
rect 1720 130 1754 548
rect 1816 130 1850 548
rect -1592 37 -1558 71
rect -1172 37 -1138 71
rect -752 37 -718 71
rect -332 37 -298 71
rect 88 37 122 71
rect 508 37 542 71
rect 928 37 962 71
rect 1348 37 1382 71
rect 1768 37 1802 71
rect -1592 -71 -1558 -37
rect -1172 -71 -1138 -37
rect -752 -71 -718 -37
rect -332 -71 -298 -37
rect 88 -71 122 -37
rect 508 -71 542 -37
rect 928 -71 962 -37
rect 1348 -71 1382 -37
rect 1768 -71 1802 -37
rect -1850 -548 -1816 -130
rect -1754 -548 -1720 -130
rect -1640 -548 -1606 -130
rect -1544 -548 -1510 -130
rect -1430 -548 -1396 -130
rect -1334 -548 -1300 -130
rect -1220 -548 -1186 -130
rect -1124 -548 -1090 -130
rect -1010 -548 -976 -130
rect -914 -548 -880 -130
rect -800 -548 -766 -130
rect -704 -548 -670 -130
rect -590 -548 -556 -130
rect -494 -548 -460 -130
rect -380 -548 -346 -130
rect -284 -548 -250 -130
rect -170 -548 -136 -130
rect -74 -548 -40 -130
rect 40 -548 74 -130
rect 136 -548 170 -130
rect 250 -548 284 -130
rect 346 -548 380 -130
rect 460 -548 494 -130
rect 556 -548 590 -130
rect 670 -548 704 -130
rect 766 -548 800 -130
rect 880 -548 914 -130
rect 976 -548 1010 -130
rect 1090 -548 1124 -130
rect 1186 -548 1220 -130
rect 1300 -548 1334 -130
rect 1396 -548 1430 -130
rect 1510 -548 1544 -130
rect 1606 -548 1640 -130
rect 1720 -548 1754 -130
rect 1816 -548 1850 -130
rect -1802 -641 -1768 -607
rect -1382 -641 -1348 -607
rect -962 -641 -928 -607
rect -542 -641 -508 -607
rect -122 -641 -88 -607
rect 298 -641 332 -607
rect 718 -641 752 -607
rect 1138 -641 1172 -607
rect 1558 -641 1592 -607
<< metal1 >>
rect -1814 641 -1756 647
rect -1814 607 -1802 641
rect -1768 607 -1756 641
rect -1814 601 -1756 607
rect -1394 641 -1336 647
rect -1394 607 -1382 641
rect -1348 607 -1336 641
rect -1394 601 -1336 607
rect -974 641 -916 647
rect -974 607 -962 641
rect -928 607 -916 641
rect -974 601 -916 607
rect -554 641 -496 647
rect -554 607 -542 641
rect -508 607 -496 641
rect -554 601 -496 607
rect -134 641 -76 647
rect -134 607 -122 641
rect -88 607 -76 641
rect -134 601 -76 607
rect 286 641 344 647
rect 286 607 298 641
rect 332 607 344 641
rect 286 601 344 607
rect 706 641 764 647
rect 706 607 718 641
rect 752 607 764 641
rect 706 601 764 607
rect 1126 641 1184 647
rect 1126 607 1138 641
rect 1172 607 1184 641
rect 1126 601 1184 607
rect 1546 641 1604 647
rect 1546 607 1558 641
rect 1592 607 1604 641
rect 1546 601 1604 607
rect -1856 548 -1810 560
rect -1856 130 -1850 548
rect -1816 130 -1810 548
rect -1856 118 -1810 130
rect -1760 548 -1714 560
rect -1760 130 -1754 548
rect -1720 130 -1714 548
rect -1760 118 -1714 130
rect -1646 548 -1600 560
rect -1646 130 -1640 548
rect -1606 130 -1600 548
rect -1646 118 -1600 130
rect -1550 548 -1504 560
rect -1550 130 -1544 548
rect -1510 130 -1504 548
rect -1550 118 -1504 130
rect -1436 548 -1390 560
rect -1436 130 -1430 548
rect -1396 130 -1390 548
rect -1436 118 -1390 130
rect -1340 548 -1294 560
rect -1340 130 -1334 548
rect -1300 130 -1294 548
rect -1340 118 -1294 130
rect -1226 548 -1180 560
rect -1226 130 -1220 548
rect -1186 130 -1180 548
rect -1226 118 -1180 130
rect -1130 548 -1084 560
rect -1130 130 -1124 548
rect -1090 130 -1084 548
rect -1130 118 -1084 130
rect -1016 548 -970 560
rect -1016 130 -1010 548
rect -976 130 -970 548
rect -1016 118 -970 130
rect -920 548 -874 560
rect -920 130 -914 548
rect -880 130 -874 548
rect -920 118 -874 130
rect -806 548 -760 560
rect -806 130 -800 548
rect -766 130 -760 548
rect -806 118 -760 130
rect -710 548 -664 560
rect -710 130 -704 548
rect -670 130 -664 548
rect -710 118 -664 130
rect -596 548 -550 560
rect -596 130 -590 548
rect -556 130 -550 548
rect -596 118 -550 130
rect -500 548 -454 560
rect -500 130 -494 548
rect -460 130 -454 548
rect -500 118 -454 130
rect -386 548 -340 560
rect -386 130 -380 548
rect -346 130 -340 548
rect -386 118 -340 130
rect -290 548 -244 560
rect -290 130 -284 548
rect -250 130 -244 548
rect -290 118 -244 130
rect -176 548 -130 560
rect -176 130 -170 548
rect -136 130 -130 548
rect -176 118 -130 130
rect -80 548 -34 560
rect -80 130 -74 548
rect -40 130 -34 548
rect -80 118 -34 130
rect 34 548 80 560
rect 34 130 40 548
rect 74 130 80 548
rect 34 118 80 130
rect 130 548 176 560
rect 130 130 136 548
rect 170 130 176 548
rect 130 118 176 130
rect 244 548 290 560
rect 244 130 250 548
rect 284 130 290 548
rect 244 118 290 130
rect 340 548 386 560
rect 340 130 346 548
rect 380 130 386 548
rect 340 118 386 130
rect 454 548 500 560
rect 454 130 460 548
rect 494 130 500 548
rect 454 118 500 130
rect 550 548 596 560
rect 550 130 556 548
rect 590 130 596 548
rect 550 118 596 130
rect 664 548 710 560
rect 664 130 670 548
rect 704 130 710 548
rect 664 118 710 130
rect 760 548 806 560
rect 760 130 766 548
rect 800 130 806 548
rect 760 118 806 130
rect 874 548 920 560
rect 874 130 880 548
rect 914 130 920 548
rect 874 118 920 130
rect 970 548 1016 560
rect 970 130 976 548
rect 1010 130 1016 548
rect 970 118 1016 130
rect 1084 548 1130 560
rect 1084 130 1090 548
rect 1124 130 1130 548
rect 1084 118 1130 130
rect 1180 548 1226 560
rect 1180 130 1186 548
rect 1220 130 1226 548
rect 1180 118 1226 130
rect 1294 548 1340 560
rect 1294 130 1300 548
rect 1334 130 1340 548
rect 1294 118 1340 130
rect 1390 548 1436 560
rect 1390 130 1396 548
rect 1430 130 1436 548
rect 1390 118 1436 130
rect 1504 548 1550 560
rect 1504 130 1510 548
rect 1544 130 1550 548
rect 1504 118 1550 130
rect 1600 548 1646 560
rect 1600 130 1606 548
rect 1640 130 1646 548
rect 1600 118 1646 130
rect 1714 548 1760 560
rect 1714 130 1720 548
rect 1754 130 1760 548
rect 1714 118 1760 130
rect 1810 548 1856 560
rect 1810 130 1816 548
rect 1850 130 1856 548
rect 1810 118 1856 130
rect -1604 71 -1546 77
rect -1604 37 -1592 71
rect -1558 37 -1546 71
rect -1604 31 -1546 37
rect -1184 71 -1126 77
rect -1184 37 -1172 71
rect -1138 37 -1126 71
rect -1184 31 -1126 37
rect -764 71 -706 77
rect -764 37 -752 71
rect -718 37 -706 71
rect -764 31 -706 37
rect -344 71 -286 77
rect -344 37 -332 71
rect -298 37 -286 71
rect -344 31 -286 37
rect 76 71 134 77
rect 76 37 88 71
rect 122 37 134 71
rect 76 31 134 37
rect 496 71 554 77
rect 496 37 508 71
rect 542 37 554 71
rect 496 31 554 37
rect 916 71 974 77
rect 916 37 928 71
rect 962 37 974 71
rect 916 31 974 37
rect 1336 71 1394 77
rect 1336 37 1348 71
rect 1382 37 1394 71
rect 1336 31 1394 37
rect 1756 71 1814 77
rect 1756 37 1768 71
rect 1802 37 1814 71
rect 1756 31 1814 37
rect -1604 -37 -1546 -31
rect -1604 -71 -1592 -37
rect -1558 -71 -1546 -37
rect -1604 -77 -1546 -71
rect -1184 -37 -1126 -31
rect -1184 -71 -1172 -37
rect -1138 -71 -1126 -37
rect -1184 -77 -1126 -71
rect -764 -37 -706 -31
rect -764 -71 -752 -37
rect -718 -71 -706 -37
rect -764 -77 -706 -71
rect -344 -37 -286 -31
rect -344 -71 -332 -37
rect -298 -71 -286 -37
rect -344 -77 -286 -71
rect 76 -37 134 -31
rect 76 -71 88 -37
rect 122 -71 134 -37
rect 76 -77 134 -71
rect 496 -37 554 -31
rect 496 -71 508 -37
rect 542 -71 554 -37
rect 496 -77 554 -71
rect 916 -37 974 -31
rect 916 -71 928 -37
rect 962 -71 974 -37
rect 916 -77 974 -71
rect 1336 -37 1394 -31
rect 1336 -71 1348 -37
rect 1382 -71 1394 -37
rect 1336 -77 1394 -71
rect 1756 -37 1814 -31
rect 1756 -71 1768 -37
rect 1802 -71 1814 -37
rect 1756 -77 1814 -71
rect -1856 -130 -1810 -118
rect -1856 -548 -1850 -130
rect -1816 -548 -1810 -130
rect -1856 -560 -1810 -548
rect -1760 -130 -1714 -118
rect -1760 -548 -1754 -130
rect -1720 -548 -1714 -130
rect -1760 -560 -1714 -548
rect -1646 -130 -1600 -118
rect -1646 -548 -1640 -130
rect -1606 -548 -1600 -130
rect -1646 -560 -1600 -548
rect -1550 -130 -1504 -118
rect -1550 -548 -1544 -130
rect -1510 -548 -1504 -130
rect -1550 -560 -1504 -548
rect -1436 -130 -1390 -118
rect -1436 -548 -1430 -130
rect -1396 -548 -1390 -130
rect -1436 -560 -1390 -548
rect -1340 -130 -1294 -118
rect -1340 -548 -1334 -130
rect -1300 -548 -1294 -130
rect -1340 -560 -1294 -548
rect -1226 -130 -1180 -118
rect -1226 -548 -1220 -130
rect -1186 -548 -1180 -130
rect -1226 -560 -1180 -548
rect -1130 -130 -1084 -118
rect -1130 -548 -1124 -130
rect -1090 -548 -1084 -130
rect -1130 -560 -1084 -548
rect -1016 -130 -970 -118
rect -1016 -548 -1010 -130
rect -976 -548 -970 -130
rect -1016 -560 -970 -548
rect -920 -130 -874 -118
rect -920 -548 -914 -130
rect -880 -548 -874 -130
rect -920 -560 -874 -548
rect -806 -130 -760 -118
rect -806 -548 -800 -130
rect -766 -548 -760 -130
rect -806 -560 -760 -548
rect -710 -130 -664 -118
rect -710 -548 -704 -130
rect -670 -548 -664 -130
rect -710 -560 -664 -548
rect -596 -130 -550 -118
rect -596 -548 -590 -130
rect -556 -548 -550 -130
rect -596 -560 -550 -548
rect -500 -130 -454 -118
rect -500 -548 -494 -130
rect -460 -548 -454 -130
rect -500 -560 -454 -548
rect -386 -130 -340 -118
rect -386 -548 -380 -130
rect -346 -548 -340 -130
rect -386 -560 -340 -548
rect -290 -130 -244 -118
rect -290 -548 -284 -130
rect -250 -548 -244 -130
rect -290 -560 -244 -548
rect -176 -130 -130 -118
rect -176 -548 -170 -130
rect -136 -548 -130 -130
rect -176 -560 -130 -548
rect -80 -130 -34 -118
rect -80 -548 -74 -130
rect -40 -548 -34 -130
rect -80 -560 -34 -548
rect 34 -130 80 -118
rect 34 -548 40 -130
rect 74 -548 80 -130
rect 34 -560 80 -548
rect 130 -130 176 -118
rect 130 -548 136 -130
rect 170 -548 176 -130
rect 130 -560 176 -548
rect 244 -130 290 -118
rect 244 -548 250 -130
rect 284 -548 290 -130
rect 244 -560 290 -548
rect 340 -130 386 -118
rect 340 -548 346 -130
rect 380 -548 386 -130
rect 340 -560 386 -548
rect 454 -130 500 -118
rect 454 -548 460 -130
rect 494 -548 500 -130
rect 454 -560 500 -548
rect 550 -130 596 -118
rect 550 -548 556 -130
rect 590 -548 596 -130
rect 550 -560 596 -548
rect 664 -130 710 -118
rect 664 -548 670 -130
rect 704 -548 710 -130
rect 664 -560 710 -548
rect 760 -130 806 -118
rect 760 -548 766 -130
rect 800 -548 806 -130
rect 760 -560 806 -548
rect 874 -130 920 -118
rect 874 -548 880 -130
rect 914 -548 920 -130
rect 874 -560 920 -548
rect 970 -130 1016 -118
rect 970 -548 976 -130
rect 1010 -548 1016 -130
rect 970 -560 1016 -548
rect 1084 -130 1130 -118
rect 1084 -548 1090 -130
rect 1124 -548 1130 -130
rect 1084 -560 1130 -548
rect 1180 -130 1226 -118
rect 1180 -548 1186 -130
rect 1220 -548 1226 -130
rect 1180 -560 1226 -548
rect 1294 -130 1340 -118
rect 1294 -548 1300 -130
rect 1334 -548 1340 -130
rect 1294 -560 1340 -548
rect 1390 -130 1436 -118
rect 1390 -548 1396 -130
rect 1430 -548 1436 -130
rect 1390 -560 1436 -548
rect 1504 -130 1550 -118
rect 1504 -548 1510 -130
rect 1544 -548 1550 -130
rect 1504 -560 1550 -548
rect 1600 -130 1646 -118
rect 1600 -548 1606 -130
rect 1640 -548 1646 -130
rect 1600 -560 1646 -548
rect 1714 -130 1760 -118
rect 1714 -548 1720 -130
rect 1754 -548 1760 -130
rect 1714 -560 1760 -548
rect 1810 -130 1856 -118
rect 1810 -548 1816 -130
rect 1850 -548 1856 -130
rect 1810 -560 1856 -548
rect -1814 -607 -1756 -601
rect -1814 -641 -1802 -607
rect -1768 -641 -1756 -607
rect -1814 -647 -1756 -641
rect -1394 -607 -1336 -601
rect -1394 -641 -1382 -607
rect -1348 -641 -1336 -607
rect -1394 -647 -1336 -641
rect -974 -607 -916 -601
rect -974 -641 -962 -607
rect -928 -641 -916 -607
rect -974 -647 -916 -641
rect -554 -607 -496 -601
rect -554 -641 -542 -607
rect -508 -641 -496 -607
rect -554 -647 -496 -641
rect -134 -607 -76 -601
rect -134 -641 -122 -607
rect -88 -641 -76 -607
rect -134 -647 -76 -641
rect 286 -607 344 -601
rect 286 -641 298 -607
rect 332 -641 344 -607
rect 286 -647 344 -641
rect 706 -607 764 -601
rect 706 -641 718 -607
rect 752 -641 764 -607
rect 706 -647 764 -641
rect 1126 -607 1184 -601
rect 1126 -641 1138 -607
rect 1172 -641 1184 -607
rect 1126 -647 1184 -641
rect 1546 -607 1604 -601
rect 1546 -641 1558 -607
rect 1592 -641 1604 -607
rect 1546 -647 1604 -641
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1947 -726 1947 726
string parameters w 2.21 l 0.15 m 2 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
