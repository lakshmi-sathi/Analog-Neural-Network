magic
tech sky130A
magscale 1 2
timestamp 1628059907
<< error_p >>
rect -29 1321 29 1327
rect -29 1287 -17 1321
rect -29 1281 29 1287
<< pwell >>
rect -211 -1459 211 1459
<< nmos >>
rect -15 -1311 15 1249
<< ndiff >>
rect -73 1237 -15 1249
rect -73 -1299 -61 1237
rect -27 -1299 -15 1237
rect -73 -1311 -15 -1299
rect 15 1237 73 1249
rect 15 -1299 27 1237
rect 61 -1299 73 1237
rect 15 -1311 73 -1299
<< ndiffc >>
rect -61 -1299 -27 1237
rect 27 -1299 61 1237
<< psubdiff >>
rect -175 1389 -79 1423
rect 79 1389 175 1423
rect -175 1327 -141 1389
rect 141 1327 175 1389
rect -175 -1389 -141 -1327
rect 141 -1389 175 -1327
rect -175 -1423 -79 -1389
rect 79 -1423 175 -1389
<< psubdiffcont >>
rect -79 1389 79 1423
rect -175 -1327 -141 1327
rect 141 -1327 175 1327
rect -79 -1423 79 -1389
<< poly >>
rect -33 1321 33 1337
rect -33 1287 -17 1321
rect 17 1287 33 1321
rect -33 1271 33 1287
rect -15 1249 15 1271
rect -15 -1337 15 -1311
<< polycont >>
rect -17 1287 17 1321
<< locali >>
rect -175 1389 -79 1423
rect 79 1389 175 1423
rect -175 1327 -141 1389
rect 141 1327 175 1389
rect -33 1287 -17 1321
rect 17 1287 33 1321
rect -61 1237 -27 1253
rect -61 -1315 -27 -1299
rect 27 1237 61 1253
rect 27 -1315 61 -1299
rect -175 -1389 -141 -1327
rect 141 -1389 175 -1327
rect -175 -1423 -79 -1389
rect 79 -1423 175 -1389
<< viali >>
rect -17 1287 17 1321
rect -61 -1299 -27 1237
rect 27 -1299 61 1237
<< metal1 >>
rect -29 1321 29 1327
rect -29 1287 -17 1321
rect 17 1287 29 1321
rect -29 1281 29 1287
rect -67 1237 -21 1249
rect -67 -1299 -61 1237
rect -27 -1299 -21 1237
rect -67 -1311 -21 -1299
rect 21 1237 67 1249
rect 21 -1299 27 1237
rect 61 -1299 67 1237
rect 21 -1311 67 -1299
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -1406 158 1406
string parameters w 12.8 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
