magic
tech sky130A
magscale 1 2
timestamp 1628080314
<< poly >>
rect 1196 371 1226 429
rect 1143 367 1226 371
rect 1127 341 1226 367
rect 247 -342 277 -281
rect 247 -372 318 -342
<< viali >>
rect 464 1464 1288 1522
rect 47 -597 1691 -525
<< metal1 >>
rect 452 1522 1300 1528
rect 452 1464 464 1522
rect 1288 1464 1300 1522
rect 452 1458 1300 1464
rect 1425 1378 1548 1383
rect 606 1332 1548 1378
rect 456 938 466 1292
rect 520 938 530 1292
rect 648 938 658 1292
rect 712 938 722 1292
rect 840 938 850 1292
rect 904 938 914 1292
rect 1032 938 1042 1292
rect 1096 938 1106 1292
rect 1224 938 1234 1292
rect 1288 938 1298 1292
rect 544 442 554 782
rect 620 442 630 782
rect 736 442 746 782
rect 812 442 822 782
rect 928 442 938 782
rect 1004 442 1014 782
rect 1120 442 1130 782
rect 1196 442 1206 782
rect 1425 386 1548 1332
rect 1660 684 1952 1006
rect 506 340 1548 386
rect 324 140 334 208
rect 766 140 776 208
rect 1425 153 1548 340
rect 1425 152 1705 153
rect 334 20 762 140
rect 1425 90 1798 152
rect 974 74 1798 90
rect 974 14 1796 74
rect 1396 8 1796 14
rect 1486 6 1666 8
rect 244 -294 296 -230
rect 448 -242 458 -190
rect 776 -242 786 -190
rect 944 -340 954 -280
rect 1272 -340 1282 -280
rect 1486 -318 1574 6
rect 448 -430 458 -378
rect 776 -430 786 -378
rect 1380 -398 1574 -318
rect 41 -519 1697 -504
rect 35 -525 1703 -519
rect 35 -597 47 -525
rect 1691 -597 1703 -525
rect 35 -603 1703 -597
rect 41 -605 1697 -603
<< via1 >>
rect 464 1464 1288 1522
rect 466 938 520 1292
rect 658 938 712 1292
rect 850 938 904 1292
rect 1042 938 1096 1292
rect 1234 938 1288 1292
rect 554 442 620 782
rect 746 442 812 782
rect 938 442 1004 782
rect 1130 442 1196 782
rect 334 140 766 208
rect 458 -242 776 -190
rect 954 -340 1272 -280
rect 458 -430 776 -378
rect 47 -597 1691 -525
<< metal2 >>
rect -52 1558 1820 1584
rect -54 1522 1824 1558
rect -54 1478 464 1522
rect 462 1464 464 1478
rect 1288 1478 1824 1522
rect 1288 1464 1296 1478
rect 462 1446 1296 1464
rect 464 1408 1296 1446
rect 462 1292 1296 1408
rect 462 938 466 1292
rect 520 938 658 1292
rect 712 938 850 1292
rect 904 938 1042 1292
rect 1096 938 1234 1292
rect 1288 1220 1296 1292
rect 1288 938 1290 1220
rect 462 934 1290 938
rect 466 928 520 934
rect 658 928 712 934
rect 850 928 904 934
rect 1042 928 1096 934
rect 1234 928 1288 934
rect 554 782 620 792
rect 554 432 620 442
rect 746 782 812 792
rect 746 432 812 442
rect 938 782 1004 792
rect 938 432 1004 442
rect 1130 782 1196 792
rect 1130 432 1196 442
rect 334 208 766 218
rect 334 130 766 140
rect 460 -180 776 -178
rect 458 -190 776 -180
rect 458 -252 776 -242
rect 460 -368 776 -252
rect 954 -280 1272 -270
rect 954 -350 1272 -340
rect 458 -378 776 -368
rect 458 -440 776 -430
rect 460 -515 776 -440
rect 47 -525 1691 -515
rect -63 -597 47 -583
rect 1691 -597 1811 -583
rect -63 -721 1811 -597
<< via2 >>
rect 554 442 620 782
rect 746 442 812 782
rect 938 442 1004 782
rect 1130 442 1196 782
rect 334 140 766 208
rect 954 -340 1272 -280
<< metal3 >>
rect 544 784 630 787
rect 736 784 822 787
rect 928 784 1014 787
rect 1120 784 1206 787
rect 538 782 1210 784
rect 538 442 554 782
rect 620 442 746 782
rect 812 442 938 782
rect 1004 442 1130 782
rect 1196 442 1210 782
rect 538 226 1210 442
rect 30 208 1210 226
rect 30 140 334 208
rect 766 140 1210 208
rect 30 138 1210 140
rect 35 136 1210 138
rect 324 135 776 136
rect 954 -275 1210 136
rect 944 -280 1282 -275
rect 944 -340 954 -280
rect 1272 -340 1282 -280
rect 944 -345 1282 -340
rect 954 -346 1210 -345
use sky130_fd_pr__nfet_01v8_XG2GE7  sky130_fd_pr__nfet_01v8_XG2GE7_0
timestamp 1628080314
transform 0 1 838 -1 0 -309
box -263 -720 263 720
use sky130_fd_pr__pfet_01v8_396TWK  sky130_fd_pr__pfet_01v8_396TWK_0
timestamp 1628080314
transform 1 0 875 0 1 859
box -551 -649 551 649
use sky130_fd_pr__res_high_po_0p35_C72MAQ  sky130_fd_pr__res_high_po_0p35_C72MAQ_0
timestamp 1628058135
transform 0 1 864 -1 0 53
box -37 -532 37 532
use sky130_fd_pr__res_high_po_0p69_7JPRER  sky130_fd_pr__res_high_po_0p69_7JPRER_0
timestamp 1628069922
transform 1 0 1719 0 1 543
box -71 -527 71 527
<< labels >>
rlabel metal2 -63 -721 1811 -597 1 GND
port 2 n
rlabel metal3 38 142 182 222 1 Out
port 6 n
rlabel metal1 1810 692 1948 1002 1 In
port 5 n
rlabel metal2 -52 1480 1818 1584 1 VDD
port 1 n
<< end >>
