magic
tech sky130A
magscale 1 2
timestamp 1627800606
<< nwell >>
rect -24 -640 4314 -636
rect -52 -1438 4314 -640
rect -52 -1442 348 -1438
<< psubdiff >>
rect 252 -1706 276 -1502
rect 2286 -1706 2310 -1502
<< nsubdiff >>
rect -16 -706 32 -682
rect 30 -1366 32 -706
rect 4230 -702 4278 -678
rect -16 -1390 32 -1366
rect 4276 -1362 4278 -702
rect 4230 -1386 4278 -1362
<< psubdiffcont >>
rect 276 -1706 2286 -1502
<< nsubdiffcont >>
rect -16 -1366 30 -706
rect 4230 -1362 4276 -702
<< poly >>
rect 4084 -1393 4114 -1341
rect 4027 -1423 4114 -1393
<< locali >>
rect 88 -544 4166 -538
rect 88 -592 96 -544
rect 4160 -592 4166 -544
rect 88 -600 4166 -592
rect -16 -706 32 -682
rect 30 -1366 32 -706
rect -16 -1390 32 -1366
rect 4230 -702 4278 -678
rect 4276 -1362 4278 -702
rect 4230 -1386 4278 -1362
rect 260 -1706 276 -1502
rect 2286 -1706 2302 -1502
<< viali >>
rect 96 -592 4160 -544
<< metal1 >>
rect 84 -594 96 -538
rect 4160 -594 4172 -538
rect 84 -604 4172 -594
rect 226 -650 4130 -642
rect 226 -704 4132 -650
rect 226 -706 4130 -704
rect 82 -1032 88 -742
rect 144 -1032 150 -742
rect 274 -1032 280 -742
rect 336 -1032 342 -742
rect 466 -1032 472 -742
rect 528 -1032 534 -742
rect 658 -1032 664 -742
rect 720 -1032 726 -742
rect 850 -1032 856 -742
rect 912 -1032 918 -742
rect 1042 -1032 1048 -742
rect 1104 -1032 1110 -742
rect 1234 -1032 1240 -742
rect 1296 -1032 1302 -742
rect 1426 -1032 1432 -742
rect 1488 -1032 1494 -742
rect 1618 -1032 1624 -742
rect 1680 -1032 1686 -742
rect 1810 -1032 1816 -742
rect 1872 -1032 1878 -742
rect 2002 -1032 2008 -742
rect 2064 -1032 2070 -742
rect 2194 -1032 2200 -742
rect 2256 -1032 2262 -742
rect 2386 -1032 2392 -742
rect 2448 -1032 2454 -742
rect 2578 -1032 2584 -742
rect 2640 -1032 2646 -742
rect 2770 -1032 2776 -742
rect 2832 -1032 2838 -742
rect 2962 -1032 2968 -742
rect 3024 -1032 3030 -742
rect 3154 -1032 3160 -742
rect 3216 -1032 3222 -742
rect 3346 -1032 3352 -742
rect 3408 -1032 3414 -742
rect 3538 -1032 3544 -742
rect 3600 -1032 3606 -742
rect 3730 -1032 3736 -742
rect 3792 -1032 3798 -742
rect 3922 -1032 3928 -742
rect 3984 -1032 3990 -742
rect 4114 -1032 4120 -742
rect 4176 -1032 4182 -742
rect 180 -1342 186 -1080
rect 238 -1342 244 -1080
rect 180 -1350 244 -1342
rect 372 -1342 378 -1080
rect 430 -1342 436 -1080
rect 372 -1350 436 -1342
rect 564 -1342 570 -1080
rect 622 -1342 628 -1080
rect 564 -1350 628 -1342
rect 756 -1342 762 -1080
rect 814 -1342 820 -1080
rect 756 -1350 820 -1342
rect 948 -1342 954 -1080
rect 1006 -1342 1012 -1080
rect 948 -1350 1012 -1342
rect 1140 -1342 1146 -1080
rect 1198 -1342 1204 -1080
rect 1140 -1350 1204 -1342
rect 1332 -1342 1338 -1080
rect 1390 -1342 1396 -1080
rect 1332 -1350 1396 -1342
rect 1524 -1342 1530 -1080
rect 1582 -1342 1588 -1080
rect 1524 -1350 1588 -1342
rect 1716 -1342 1722 -1080
rect 1774 -1342 1780 -1080
rect 1716 -1350 1780 -1342
rect 1908 -1342 1914 -1080
rect 1966 -1342 1972 -1080
rect 1908 -1350 1972 -1342
rect 2100 -1342 2106 -1080
rect 2158 -1342 2164 -1080
rect 2100 -1350 2164 -1342
rect 2292 -1342 2298 -1080
rect 2350 -1342 2356 -1080
rect 2292 -1350 2356 -1342
rect 2484 -1342 2490 -1080
rect 2542 -1342 2548 -1080
rect 2484 -1350 2548 -1342
rect 2676 -1342 2682 -1080
rect 2734 -1342 2740 -1080
rect 2676 -1350 2740 -1342
rect 2868 -1342 2874 -1080
rect 2926 -1342 2932 -1080
rect 2868 -1350 2932 -1342
rect 3060 -1342 3066 -1080
rect 3118 -1342 3124 -1080
rect 3060 -1350 3124 -1342
rect 3252 -1342 3258 -1080
rect 3310 -1342 3316 -1080
rect 3252 -1350 3316 -1342
rect 3444 -1342 3450 -1080
rect 3502 -1342 3508 -1080
rect 3444 -1350 3508 -1342
rect 3636 -1342 3642 -1080
rect 3694 -1342 3700 -1080
rect 3636 -1350 3700 -1342
rect 3828 -1342 3834 -1080
rect 3886 -1342 3892 -1080
rect 3828 -1350 3892 -1342
rect 4020 -1342 4026 -1080
rect 4078 -1342 4084 -1080
rect 4020 -1350 4084 -1342
rect 132 -1432 4036 -1378
<< via1 >>
rect 96 -544 4160 -538
rect 96 -592 4160 -544
rect 96 -594 4160 -592
rect 88 -1032 144 -742
rect 280 -1032 336 -742
rect 472 -1032 528 -742
rect 664 -1032 720 -742
rect 856 -1032 912 -742
rect 1048 -1032 1104 -742
rect 1240 -1032 1296 -742
rect 1432 -1032 1488 -742
rect 1624 -1032 1680 -742
rect 1816 -1032 1872 -742
rect 2008 -1032 2064 -742
rect 2200 -1032 2256 -742
rect 2392 -1032 2448 -742
rect 2584 -1032 2640 -742
rect 2776 -1032 2832 -742
rect 2968 -1032 3024 -742
rect 3160 -1032 3216 -742
rect 3352 -1032 3408 -742
rect 3544 -1032 3600 -742
rect 3736 -1032 3792 -742
rect 3928 -1032 3984 -742
rect 4120 -1032 4176 -742
rect 186 -1342 238 -1080
rect 378 -1342 430 -1080
rect 570 -1342 622 -1080
rect 762 -1342 814 -1080
rect 954 -1342 1006 -1080
rect 1146 -1342 1198 -1080
rect 1338 -1342 1390 -1080
rect 1530 -1342 1582 -1080
rect 1722 -1342 1774 -1080
rect 1914 -1342 1966 -1080
rect 2106 -1342 2158 -1080
rect 2298 -1342 2350 -1080
rect 2490 -1342 2542 -1080
rect 2682 -1342 2734 -1080
rect 2874 -1342 2926 -1080
rect 3066 -1342 3118 -1080
rect 3258 -1342 3310 -1080
rect 3450 -1342 3502 -1080
rect 3642 -1342 3694 -1080
rect 3834 -1342 3886 -1080
rect 4026 -1342 4078 -1080
<< metal2 >>
rect 82 -538 4182 -516
rect 82 -594 96 -538
rect 4160 -594 4182 -538
rect 82 -622 4182 -594
rect 82 -742 150 -622
rect 82 -1032 88 -742
rect 144 -1032 150 -742
rect 274 -742 342 -622
rect 274 -1032 280 -742
rect 336 -1032 342 -742
rect 466 -742 534 -622
rect 466 -1032 472 -742
rect 528 -1032 534 -742
rect 658 -742 726 -622
rect 658 -1032 664 -742
rect 720 -1032 726 -742
rect 850 -742 918 -622
rect 850 -1032 856 -742
rect 912 -1032 918 -742
rect 1042 -742 1110 -622
rect 1042 -1032 1048 -742
rect 1104 -1032 1110 -742
rect 1234 -742 1302 -622
rect 1234 -1032 1240 -742
rect 1296 -1032 1302 -742
rect 1426 -742 1494 -622
rect 1426 -1032 1432 -742
rect 1488 -1032 1494 -742
rect 1618 -742 1686 -622
rect 1618 -1032 1624 -742
rect 1680 -1032 1686 -742
rect 1810 -742 1878 -622
rect 1810 -1032 1816 -742
rect 1872 -1032 1878 -742
rect 2002 -742 2070 -622
rect 2002 -1032 2008 -742
rect 2064 -1032 2070 -742
rect 2194 -742 2262 -622
rect 2194 -1032 2200 -742
rect 2256 -1032 2262 -742
rect 2386 -742 2454 -622
rect 2386 -1032 2392 -742
rect 2448 -1032 2454 -742
rect 2578 -742 2646 -622
rect 2578 -1032 2584 -742
rect 2640 -1032 2646 -742
rect 2770 -742 2838 -622
rect 2770 -1032 2776 -742
rect 2832 -1032 2838 -742
rect 2962 -742 3030 -622
rect 2962 -1032 2968 -742
rect 3024 -1032 3030 -742
rect 3154 -742 3222 -622
rect 3154 -1032 3160 -742
rect 3216 -1032 3222 -742
rect 3346 -742 3414 -622
rect 3346 -1032 3352 -742
rect 3408 -1032 3414 -742
rect 3538 -742 3606 -622
rect 3538 -1032 3544 -742
rect 3600 -1032 3606 -742
rect 3730 -742 3798 -622
rect 3730 -1032 3736 -742
rect 3792 -1032 3798 -742
rect 3922 -742 3990 -622
rect 3922 -1032 3928 -742
rect 3984 -1032 3990 -742
rect 4114 -742 4182 -622
rect 4114 -1032 4120 -742
rect 4176 -1032 4182 -742
rect 180 -1080 244 -1070
rect 180 -1340 184 -1080
rect 240 -1340 244 -1080
rect 180 -1342 186 -1340
rect 238 -1342 244 -1340
rect 180 -1350 244 -1342
rect 372 -1080 436 -1070
rect 372 -1340 376 -1080
rect 432 -1340 436 -1080
rect 372 -1342 378 -1340
rect 430 -1342 436 -1340
rect 372 -1350 436 -1342
rect 564 -1080 628 -1070
rect 564 -1340 568 -1080
rect 624 -1340 628 -1080
rect 564 -1342 570 -1340
rect 622 -1342 628 -1340
rect 564 -1350 628 -1342
rect 756 -1080 820 -1070
rect 756 -1340 760 -1080
rect 816 -1340 820 -1080
rect 756 -1342 762 -1340
rect 814 -1342 820 -1340
rect 756 -1350 820 -1342
rect 948 -1080 1012 -1070
rect 948 -1340 952 -1080
rect 1008 -1340 1012 -1080
rect 948 -1342 954 -1340
rect 1006 -1342 1012 -1340
rect 948 -1350 1012 -1342
rect 1140 -1080 1204 -1070
rect 1140 -1340 1144 -1080
rect 1200 -1340 1204 -1080
rect 1140 -1342 1146 -1340
rect 1198 -1342 1204 -1340
rect 1140 -1350 1204 -1342
rect 1332 -1080 1396 -1070
rect 1332 -1340 1336 -1080
rect 1392 -1340 1396 -1080
rect 1332 -1342 1338 -1340
rect 1390 -1342 1396 -1340
rect 1332 -1350 1396 -1342
rect 1524 -1080 1588 -1070
rect 1524 -1340 1528 -1080
rect 1584 -1340 1588 -1080
rect 1524 -1342 1530 -1340
rect 1582 -1342 1588 -1340
rect 1524 -1350 1588 -1342
rect 1716 -1080 1780 -1070
rect 1716 -1340 1720 -1080
rect 1776 -1340 1780 -1080
rect 1716 -1342 1722 -1340
rect 1774 -1342 1780 -1340
rect 1716 -1350 1780 -1342
rect 1908 -1080 1972 -1070
rect 1908 -1340 1912 -1080
rect 1968 -1340 1972 -1080
rect 1908 -1342 1914 -1340
rect 1966 -1342 1972 -1340
rect 1908 -1350 1972 -1342
rect 2100 -1080 2164 -1070
rect 2100 -1340 2104 -1080
rect 2160 -1340 2164 -1080
rect 2100 -1342 2106 -1340
rect 2158 -1342 2164 -1340
rect 2100 -1350 2164 -1342
rect 2292 -1080 2356 -1070
rect 2292 -1340 2296 -1080
rect 2352 -1340 2356 -1080
rect 2292 -1342 2298 -1340
rect 2350 -1342 2356 -1340
rect 2292 -1350 2356 -1342
rect 2484 -1080 2548 -1070
rect 2484 -1340 2488 -1080
rect 2544 -1340 2548 -1080
rect 2484 -1342 2490 -1340
rect 2542 -1342 2548 -1340
rect 2484 -1350 2548 -1342
rect 2676 -1080 2740 -1070
rect 2676 -1340 2680 -1080
rect 2736 -1340 2740 -1080
rect 2676 -1342 2682 -1340
rect 2734 -1342 2740 -1340
rect 2676 -1350 2740 -1342
rect 2868 -1080 2932 -1070
rect 2868 -1340 2872 -1080
rect 2928 -1340 2932 -1080
rect 2868 -1342 2874 -1340
rect 2926 -1342 2932 -1340
rect 2868 -1350 2932 -1342
rect 3060 -1080 3124 -1070
rect 3060 -1340 3064 -1080
rect 3120 -1340 3124 -1080
rect 3060 -1342 3066 -1340
rect 3118 -1342 3124 -1340
rect 3060 -1350 3124 -1342
rect 3252 -1080 3316 -1070
rect 3252 -1340 3256 -1080
rect 3312 -1340 3316 -1080
rect 3252 -1342 3258 -1340
rect 3310 -1342 3316 -1340
rect 3252 -1350 3316 -1342
rect 3444 -1080 3508 -1070
rect 3444 -1340 3448 -1080
rect 3504 -1340 3508 -1080
rect 3444 -1342 3450 -1340
rect 3502 -1342 3508 -1340
rect 3444 -1350 3508 -1342
rect 3636 -1080 3700 -1070
rect 3636 -1340 3640 -1080
rect 3696 -1340 3700 -1080
rect 3636 -1342 3642 -1340
rect 3694 -1342 3700 -1340
rect 3636 -1350 3700 -1342
rect 3828 -1080 3892 -1070
rect 3828 -1340 3832 -1080
rect 3888 -1340 3892 -1080
rect 3828 -1342 3834 -1340
rect 3886 -1342 3892 -1340
rect 3828 -1350 3892 -1342
rect 4020 -1080 4084 -1070
rect 4020 -1340 4024 -1080
rect 4080 -1340 4084 -1080
rect 4020 -1342 4026 -1340
rect 4078 -1342 4084 -1340
rect 4020 -1350 4084 -1342
<< via2 >>
rect 184 -1340 186 -1080
rect 186 -1340 238 -1080
rect 238 -1340 240 -1080
rect 376 -1340 378 -1080
rect 378 -1340 430 -1080
rect 430 -1340 432 -1080
rect 568 -1340 570 -1080
rect 570 -1340 622 -1080
rect 622 -1340 624 -1080
rect 760 -1340 762 -1080
rect 762 -1340 814 -1080
rect 814 -1340 816 -1080
rect 952 -1340 954 -1080
rect 954 -1340 1006 -1080
rect 1006 -1340 1008 -1080
rect 1144 -1340 1146 -1080
rect 1146 -1340 1198 -1080
rect 1198 -1340 1200 -1080
rect 1336 -1340 1338 -1080
rect 1338 -1340 1390 -1080
rect 1390 -1340 1392 -1080
rect 1528 -1340 1530 -1080
rect 1530 -1340 1582 -1080
rect 1582 -1340 1584 -1080
rect 1720 -1340 1722 -1080
rect 1722 -1340 1774 -1080
rect 1774 -1340 1776 -1080
rect 1912 -1340 1914 -1080
rect 1914 -1340 1966 -1080
rect 1966 -1340 1968 -1080
rect 2104 -1340 2106 -1080
rect 2106 -1340 2158 -1080
rect 2158 -1340 2160 -1080
rect 2296 -1340 2298 -1080
rect 2298 -1340 2350 -1080
rect 2350 -1340 2352 -1080
rect 2488 -1340 2490 -1080
rect 2490 -1340 2542 -1080
rect 2542 -1340 2544 -1080
rect 2680 -1340 2682 -1080
rect 2682 -1340 2734 -1080
rect 2734 -1340 2736 -1080
rect 2872 -1340 2874 -1080
rect 2874 -1340 2926 -1080
rect 2926 -1340 2928 -1080
rect 3064 -1340 3066 -1080
rect 3066 -1340 3118 -1080
rect 3118 -1340 3120 -1080
rect 3256 -1340 3258 -1080
rect 3258 -1340 3310 -1080
rect 3310 -1340 3312 -1080
rect 3448 -1340 3450 -1080
rect 3450 -1340 3502 -1080
rect 3502 -1340 3504 -1080
rect 3640 -1340 3642 -1080
rect 3642 -1340 3694 -1080
rect 3694 -1340 3696 -1080
rect 3832 -1340 3834 -1080
rect 3834 -1340 3886 -1080
rect 3886 -1340 3888 -1080
rect 4024 -1340 4026 -1080
rect 4026 -1340 4078 -1080
rect 4078 -1340 4080 -1080
<< metal3 >>
rect 178 -1080 246 -1070
rect 178 -1340 184 -1080
rect 240 -1340 246 -1080
rect 178 -1396 246 -1340
rect 370 -1080 438 -1070
rect 370 -1340 376 -1080
rect 432 -1340 438 -1080
rect 370 -1396 438 -1340
rect 562 -1080 630 -1070
rect 562 -1340 568 -1080
rect 624 -1340 630 -1080
rect 562 -1396 630 -1340
rect 754 -1080 822 -1070
rect 754 -1340 760 -1080
rect 816 -1340 822 -1080
rect 754 -1396 822 -1340
rect 946 -1080 1014 -1070
rect 946 -1340 952 -1080
rect 1008 -1340 1014 -1080
rect 946 -1396 1014 -1340
rect 1138 -1080 1206 -1070
rect 1138 -1340 1144 -1080
rect 1200 -1340 1206 -1080
rect 1138 -1396 1206 -1340
rect 1330 -1080 1398 -1070
rect 1330 -1340 1336 -1080
rect 1392 -1340 1398 -1080
rect 1330 -1396 1398 -1340
rect 1522 -1080 1590 -1070
rect 1522 -1340 1528 -1080
rect 1584 -1340 1590 -1080
rect 1522 -1396 1590 -1340
rect 1714 -1080 1782 -1070
rect 1714 -1340 1720 -1080
rect 1776 -1340 1782 -1080
rect 1714 -1396 1782 -1340
rect 1906 -1080 1974 -1072
rect 1906 -1340 1912 -1080
rect 1968 -1340 1974 -1080
rect 1906 -1396 1974 -1340
rect 2098 -1080 2166 -1070
rect 2098 -1340 2104 -1080
rect 2160 -1340 2166 -1080
rect 2098 -1396 2166 -1340
rect 2290 -1080 2358 -1070
rect 2290 -1340 2296 -1080
rect 2352 -1340 2358 -1080
rect 2290 -1396 2358 -1340
rect 2482 -1080 2550 -1072
rect 2482 -1340 2488 -1080
rect 2544 -1340 2550 -1080
rect 2482 -1396 2550 -1340
rect 2674 -1080 2742 -1070
rect 2674 -1340 2680 -1080
rect 2736 -1340 2742 -1080
rect 2674 -1396 2742 -1340
rect 2866 -1080 2934 -1072
rect 2866 -1340 2872 -1080
rect 2928 -1340 2934 -1080
rect 2866 -1396 2934 -1340
rect 3058 -1080 3126 -1070
rect 3058 -1340 3064 -1080
rect 3120 -1340 3126 -1080
rect 3058 -1396 3126 -1340
rect 3250 -1080 3318 -1070
rect 3250 -1340 3256 -1080
rect 3312 -1340 3318 -1080
rect 3250 -1396 3318 -1340
rect 3442 -1080 3510 -1070
rect 3442 -1340 3448 -1080
rect 3504 -1340 3510 -1080
rect 3442 -1396 3510 -1340
rect 3634 -1080 3702 -1070
rect 3634 -1340 3640 -1080
rect 3696 -1340 3702 -1080
rect 3634 -1396 3702 -1340
rect 3826 -1080 3894 -1070
rect 3826 -1340 3832 -1080
rect 3888 -1340 3894 -1080
rect 3826 -1396 3894 -1340
rect 4018 -1080 4086 -1070
rect 4018 -1340 4024 -1080
rect 4080 -1340 4086 -1080
rect 4018 -1396 4086 -1340
rect 178 -1450 4088 -1396
rect 78 -1640 4180 -1450
use sky130_fd_pr__pfet_01v8_CC7KEW  sky130_fd_pr__pfet_01v8_CC7KEW_0
timestamp 1627668659
transform 1 0 2131 0 1 -1038
box -2081 -400 2081 400
<< labels >>
rlabel metal3 82 -1636 4176 -1558 1 vh
port 4 n
rlabel metal1 134 -1430 4034 -1378 1 gate
port 6 n
rlabel metal2 90 -612 4174 -524 1 VDD
port 7 n
rlabel psubdiffcont 276 -1706 2286 -1502 1 GND
<< end >>
