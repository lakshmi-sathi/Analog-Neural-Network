magic
tech sky130A
magscale 1 2
timestamp 1628056522
<< nmos >>
rect -15 -840 15 840
<< ndiff >>
rect -73 828 -15 840
rect -73 -828 -61 828
rect -27 -828 -15 828
rect -73 -840 -15 -828
rect 15 828 73 840
rect 15 -828 27 828
rect 61 -828 73 828
rect 15 -840 73 -828
<< ndiffc >>
rect -61 -828 -27 828
rect 27 -828 61 828
<< poly >>
rect -15 840 15 866
rect -15 -866 15 -840
<< locali >>
rect -61 828 -27 844
rect -61 -844 -27 -828
rect 27 828 61 844
rect 27 -844 61 -828
<< viali >>
rect -61 -828 -27 828
rect 27 -828 61 828
<< metal1 >>
rect -67 828 -21 840
rect -67 -828 -61 828
rect -27 -828 -21 828
rect -67 -840 -21 -828
rect 21 828 67 840
rect 21 -828 27 828
rect 61 -828 67 828
rect 21 -840 67 -828
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 8.4 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
