magic
tech sky130A
magscale 1 2
timestamp 1627890010
<< locali >>
rect 14006 -1292 14420 -1200
rect 14014 -2542 14428 -2450
rect 13992 -3810 14406 -3718
<< metal1 >>
rect 586 2556 1016 2578
rect 582 2072 592 2556
rect 994 2072 1016 2556
rect 586 1944 1016 2072
rect -514 1402 1016 1944
rect 586 1184 1016 1402
rect 11922 1672 12160 1674
rect 11922 1086 12374 1672
rect 12114 -1102 12374 1086
rect 13838 1550 15688 1910
rect 13838 -328 14198 1550
rect 15328 1208 15688 1550
rect 26632 1202 27262 1208
rect 26632 956 26652 1202
rect 27246 956 27262 1202
rect 26632 950 27262 956
rect 13838 -688 18768 -328
rect 614 -1498 956 -1222
rect -540 -2040 956 -1498
rect 11890 -1692 12374 -1102
rect 614 -2226 956 -2040
rect 614 -2590 626 -2226
rect 956 -2590 966 -2226
rect 614 -2604 956 -2590
rect 12114 -2942 12374 -1692
rect 14834 -1569 15196 -1565
rect 18370 -1566 18730 -688
rect 14834 -1779 14844 -1569
rect 14962 -1779 15196 -1569
rect 14834 -1787 15196 -1779
rect 18270 -1788 18730 -1566
rect 18298 -1790 18730 -1788
rect 18370 -2768 18730 -1790
rect 14840 -2818 15210 -2810
rect 12114 -2964 13044 -2942
rect 12114 -3656 12478 -2964
rect 13018 -3108 13044 -2964
rect 14836 -3012 14846 -2818
rect 14972 -3012 15210 -2818
rect 18270 -2990 18730 -2768
rect 14840 -3022 15210 -3012
rect 13018 -3336 13040 -3108
rect 13018 -3656 13044 -3336
rect 12114 -3668 13044 -3656
rect 600 -3836 926 -3830
rect 600 -4186 616 -3836
rect 914 -4186 926 -3836
rect 600 -4306 926 -4186
rect -548 -4848 936 -4306
rect 12114 -4584 12374 -3668
rect 18370 -4048 18730 -2990
rect 20194 -3860 20212 -2768
rect 20534 -3860 20552 -2768
rect 20194 -3888 20552 -3860
rect 14828 -4084 15202 -4078
rect 14818 -4280 14828 -4084
rect 14948 -4280 15202 -4084
rect 18272 -4266 18730 -4048
rect 18370 -4284 18730 -4266
rect 600 -5180 926 -4848
rect 11944 -5132 12374 -4584
rect 12114 -5136 12374 -5132
<< via1 >>
rect 592 2072 994 2556
rect 26652 956 27246 1202
rect 626 -2590 956 -2226
rect 14844 -1779 14962 -1569
rect 12478 -3656 13018 -2964
rect 14846 -3012 14972 -2818
rect 616 -4186 914 -3836
rect 20212 -3860 20534 -2768
rect 14828 -4280 14948 -4084
<< metal2 >>
rect 376 3148 29806 3151
rect 92 3021 30028 3148
rect 92 3014 1595 3021
rect 94 -2996 350 3014
rect 26040 2967 30028 3021
rect 592 2556 994 2566
rect 592 2062 994 2072
rect 26652 1202 27246 1212
rect 26652 946 27246 956
rect 1399 48 26795 130
rect 1399 -112 19024 48
rect 21144 -112 26795 48
rect 19024 -138 21144 -128
rect 19312 -414 20022 -412
rect 29622 -414 30028 2967
rect 19312 -590 30028 -414
rect 14718 -734 30028 -590
rect 14718 -777 20022 -734
rect 14708 -859 20022 -777
rect 14708 -1402 14790 -859
rect 14828 -1569 14974 -1559
rect 14828 -1779 14844 -1569
rect 14962 -1779 14974 -1569
rect 14828 -1789 14974 -1779
rect 626 -2226 956 -2216
rect 17121 -2313 17203 -859
rect 626 -2600 956 -2590
rect 14711 -2395 17203 -2313
rect 14711 -2649 14793 -2395
rect 14846 -2810 14972 -2808
rect 14838 -2818 14984 -2810
rect 12460 -2964 13056 -2940
rect 94 -3252 11994 -2996
rect 12460 -3108 12478 -2964
rect 12462 -3336 12478 -3108
rect 12460 -3656 12478 -3336
rect 13018 -3656 13056 -2964
rect 14838 -3012 14846 -2818
rect 14972 -3012 14984 -2818
rect 14838 -3020 14984 -3012
rect 14846 -3022 14972 -3020
rect 18659 -3507 18741 -859
rect 19312 -866 20022 -859
rect 20212 -2768 20534 -2758
rect 12460 -3670 13056 -3656
rect 616 -3836 914 -3826
rect 12473 -4032 13056 -3670
rect 14689 -3589 18741 -3507
rect 14689 -3925 14771 -3589
rect 19212 -3670 20212 -2940
rect 616 -4196 914 -4186
rect 12472 -4304 13056 -4032
rect 14828 -4080 14948 -4074
rect 14820 -4084 14958 -4080
rect 14820 -4280 14828 -4084
rect 14948 -4280 14958 -4084
rect 14820 -4284 14958 -4280
rect 14828 -4290 14948 -4284
rect 12473 -4900 13056 -4304
rect 12473 -5148 13048 -4900
rect 19212 -5148 19815 -3670
rect 20534 -2954 27437 -2940
rect 20534 -3658 26722 -2954
rect 27420 -3658 27437 -2954
rect 20534 -3670 27437 -3658
rect 20212 -3870 20534 -3860
rect 12473 -5697 19815 -5148
rect 19218 -5976 19910 -5966
rect 19212 -6092 19218 -6000
rect 1616 -6240 19218 -6092
rect 27612 -6000 28408 -5822
rect 19910 -6092 28408 -6000
rect 19910 -6240 28431 -6092
rect 1616 -6266 28431 -6240
<< via2 >>
rect 592 2072 994 2556
rect 26942 956 27246 1202
rect 19024 -128 21144 48
rect 626 -2590 956 -2226
rect 616 -4186 914 -3836
rect 20212 -3860 20534 -2768
rect 26722 -3658 27420 -2954
rect 19218 -6240 19910 -5976
<< metal3 >>
rect 582 2556 1004 2561
rect 582 2072 592 2556
rect 994 2072 1004 2556
rect 582 2067 1004 2072
rect 26920 1202 27276 1214
rect 26920 956 26942 1202
rect 27246 956 27276 1202
rect 11868 166 13582 486
rect 11862 -474 12740 -154
rect 616 -2226 966 -2221
rect 616 -2590 626 -2226
rect 956 -2590 966 -2226
rect 616 -2595 966 -2590
rect 12420 -3008 12740 -474
rect 13262 -1468 13582 166
rect 19000 48 21164 56
rect 19000 -128 19024 48
rect 21144 -128 21164 48
rect 19000 -136 21164 -128
rect 13262 -1750 13578 -1468
rect 13262 -1756 13670 -1750
rect 13262 -1757 13774 -1756
rect 13262 -1854 13944 -1757
rect 13774 -1855 13944 -1854
rect 13614 -3008 13962 -3006
rect 12420 -3108 13962 -3008
rect 606 -3836 924 -3831
rect 606 -4186 616 -3836
rect 914 -4186 924 -3836
rect 606 -4191 924 -4186
rect 12440 -4274 12760 -4272
rect 13776 -4274 13938 -4273
rect 12440 -4367 13938 -4274
rect 12440 -4368 13780 -4367
rect 12440 -5764 12760 -4368
rect 11882 -6084 12760 -5764
rect 19218 -5971 19914 -136
rect 20202 -2768 20544 -2763
rect 20202 -3860 20212 -2768
rect 20534 -3860 20544 -2768
rect 26920 -2949 27276 956
rect 26712 -2954 27430 -2949
rect 26712 -3658 26722 -2954
rect 27420 -3658 27430 -2954
rect 26712 -3663 27430 -3658
rect 20202 -3865 20544 -3860
rect 19208 -5976 19920 -5971
rect 19208 -6240 19218 -5976
rect 19910 -6240 19920 -5976
rect 19208 -6245 19920 -6240
<< via3 >>
rect 592 2072 994 2556
rect 626 -2590 956 -2226
rect 616 -4186 914 -3836
<< metal4 >>
rect 574 2556 13176 2580
rect 574 2072 592 2556
rect 994 2196 13176 2556
rect 994 2072 1016 2196
rect 574 2054 1016 2072
rect 12792 -1472 13176 2196
rect 30232 1966 30658 2134
rect 30188 1960 30658 1966
rect 27450 1505 30658 1960
rect 27450 1185 28143 1505
rect 30188 1504 30658 1505
rect 30232 1372 30658 1504
rect 12792 -1592 13956 -1472
rect 13278 -2224 13406 -2222
rect 610 -2226 13406 -2224
rect 610 -2590 626 -2226
rect 956 -2590 13406 -2226
rect 610 -2608 13406 -2590
rect 12938 -2614 13406 -2608
rect 13100 -2704 13406 -2614
rect 13100 -2832 13960 -2704
rect 13100 -2834 13352 -2832
rect 582 -3836 12916 -3818
rect 582 -4186 616 -3836
rect 914 -4006 12916 -3836
rect 914 -4104 13934 -4006
rect 914 -4186 12916 -4104
rect 582 -4202 12916 -4186
use voltage_div  voltage_div_0 /mnt/c/Users/LENOVO/Documents/AnalogNeuralNetwork
timestamp 1627883883
transform 1 0 20412 0 1 -3066
box 0 -2992 8012 2542
use analogneuron_invopamp_re_15kfeedbck  analogneuron_invopamp_re_15kfeedbck_0
timestamp 1627836603
transform 1 0 1354 0 1 234
box -1354 -234 10724 2910
use analogneuron_invopamp_re_15kfeedbck  analogneuron_invopamp_re_15kfeedbck_1
timestamp 1627836603
transform 1 0 1348 0 -1 -216
box -1354 -234 10724 2910
use analogneuron_invopamp_re_15kfeedbck  analogneuron_invopamp_re_15kfeedbck_2
timestamp 1627836603
transform 1 0 1358 0 1 -6032
box -1354 -234 10724 2910
use analogneuron_invopamp_re_15kfeedbck_ReLU  analogneuron_invopamp_re_15kfeedbck_ReLU_0
timestamp 1627839109
transform 1 0 16082 0 1 241
box -1354 -343 13246 2910
use mux  mux_0 /mnt/c/Users/LENOVO/Documents/AnalogNeuralNetwork
timestamp 1627111729
transform 1 0 13846 0 -1 -1597
box -22 -348 1124 429
use mux  mux_1
timestamp 1627111729
transform 1 0 13854 0 -1 -2851
box -22 -348 1124 429
use mux  mux_2
timestamp 1627111729
transform 1 0 13834 0 -1 -4119
box -22 -348 1124 429
<< labels >>
rlabel metal1 15048 -1772 15184 -1574 1 r1p1
port 1 n
rlabel metal1 15068 -3012 15204 -2814 1 r2p1
port 3 n
rlabel metal1 15052 -4278 15188 -4080 1 r3p1
port 5 n
rlabel metal1 18288 -4256 18424 -4058 1 r3p2
port 6 n
rlabel metal2 1366 3026 30014 3140 1 VDD
port 7 n
rlabel metal2 1626 -6256 28406 -6126 1 GND
port 8 n
rlabel locali 13998 -3804 14394 -3730 1 m3sel
port 9 n
rlabel locali 14022 -2534 14418 -2460 1 m2sel
port 10 n
rlabel locali 14012 -1282 14408 -1208 1 m1sel
port 11 n
rlabel metal2 1414 -90 12030 118 1 GND
port 8 n
rlabel metal2 1444 -3244 11944 -3020 1 VDD
port 7 n
rlabel metal1 -492 1428 -86 1922 1 in1
port 12 n
rlabel metal1 -514 -2020 -108 -1526 1 in2
port 13 n
rlabel metal1 -516 -4822 -110 -4328 1 in3
port 14 n
rlabel metal4 30250 1384 30628 2108 1 out
port 15 n
rlabel metal2 12482 -3690 13028 -2954 1 vcm
port 16 n
<< end >>
