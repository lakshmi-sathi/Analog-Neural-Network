magic
tech sky130A
magscale 1 2
timestamp 1627921586
<< xpolycontact >>
rect -35 99 35 531
rect -35 -531 35 -99
<< xpolyres >>
rect -35 -99 35 99
<< viali >>
rect -19 116 19 513
rect -19 -513 19 -116
<< metal1 >>
rect -25 513 25 525
rect -25 116 -19 513
rect 19 116 25 513
rect -25 104 25 116
rect -25 -116 25 -104
rect -25 -513 -19 -116
rect 19 -513 25 -116
rect -25 -525 25 -513
<< res0p35 >>
rect -37 -101 37 101
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 0.99 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 6.342k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
