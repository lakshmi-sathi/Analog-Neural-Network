magic
tech sky130A
magscale 1 2
timestamp 1628375466
<< xpolycontact >>
rect -35 86 35 518
rect -35 -518 35 -86
<< xpolyres >>
rect -35 -86 35 86
<< viali >>
rect -19 103 19 500
rect -19 -500 19 -103
<< metal1 >>
rect -25 500 25 512
rect -25 103 -19 500
rect 19 103 25 500
rect -25 91 25 103
rect -25 -103 25 -91
rect -25 -500 -19 -103
rect 19 -500 25 -103
rect -25 -512 25 -500
<< res0p35 >>
rect -37 -88 37 88
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 0.86 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.023k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
