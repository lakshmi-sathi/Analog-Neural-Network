magic
tech sky130A
magscale 1 2
timestamp 1627812750
<< nwell >>
rect -373 -420 373 420
<< nsubdiff >>
rect -337 350 -241 384
rect 241 350 337 384
rect -337 288 -303 350
rect 303 288 337 350
rect -337 -350 -303 -288
rect 303 -350 337 -288
rect -337 -384 -241 -350
rect 241 -384 337 -350
<< nsubdiffcont >>
rect -241 350 241 384
rect -337 -288 -303 288
rect 303 -288 337 288
rect -241 -384 241 -350
<< poly >>
rect -207 -203 -135 -180
rect -207 -237 -191 -203
rect -151 -237 -135 -203
rect -207 -253 -135 -237
rect 135 -203 207 -180
rect 135 -237 151 -203
rect 191 -237 207 -203
rect 135 -253 207 -237
<< polycont >>
rect -191 -237 -151 -203
rect 151 -237 191 -203
<< npolyres >>
rect -207 182 -21 254
rect -207 -180 -135 182
rect -93 -4 -21 182
rect 21 182 207 254
rect 21 -4 93 182
rect -93 -76 93 -4
rect 135 -180 207 182
<< locali >>
rect -337 350 -241 384
rect 241 350 337 384
rect -337 288 -303 350
rect 303 288 337 350
rect -207 -237 -191 -203
rect -151 -237 -135 -203
rect 135 -237 151 -203
rect 191 -237 207 -203
rect -337 -350 -303 -288
rect 303 -350 337 -288
rect -337 -384 -241 -350
rect 241 -384 337 -350
<< properties >>
string gencell sky130_fd_pr__res_generic_po
string FIXED_BBOX -320 -367 320 367
string parameters w 0.36 l 1.650 m 1 nx 4 wmin 0.330 lmin 1.650 rho 48.2 val 1.188k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 1 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
