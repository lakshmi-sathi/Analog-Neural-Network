magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< pwell >>
rect 408 -272 8000 -228
<< psubdiff >>
rect 408 -233 8000 -228
rect 408 -267 447 -233
rect 481 -267 515 -233
rect 549 -267 583 -233
rect 617 -267 651 -233
rect 685 -267 719 -233
rect 753 -267 787 -233
rect 821 -267 855 -233
rect 889 -267 923 -233
rect 957 -267 991 -233
rect 1025 -267 1059 -233
rect 1093 -267 1127 -233
rect 1161 -267 1195 -233
rect 1229 -267 1263 -233
rect 1297 -267 1331 -233
rect 1365 -267 1399 -233
rect 1433 -267 1467 -233
rect 1501 -267 1535 -233
rect 1569 -267 1603 -233
rect 1637 -267 1671 -233
rect 1705 -267 1739 -233
rect 1773 -267 1807 -233
rect 1841 -267 1875 -233
rect 1909 -267 1943 -233
rect 1977 -267 2011 -233
rect 2045 -267 2079 -233
rect 2113 -267 2147 -233
rect 2181 -267 2215 -233
rect 2249 -267 2283 -233
rect 2317 -267 2351 -233
rect 2385 -267 2419 -233
rect 2453 -267 2487 -233
rect 2521 -267 2555 -233
rect 2589 -267 2623 -233
rect 2657 -267 2691 -233
rect 2725 -267 2759 -233
rect 2793 -267 2827 -233
rect 2861 -267 2895 -233
rect 2929 -267 2963 -233
rect 2997 -267 3031 -233
rect 3065 -267 3099 -233
rect 3133 -267 3167 -233
rect 3201 -267 3235 -233
rect 3269 -267 3303 -233
rect 3337 -267 3371 -233
rect 3405 -267 3439 -233
rect 3473 -267 3507 -233
rect 3541 -267 3575 -233
rect 3609 -267 3643 -233
rect 3677 -267 3711 -233
rect 3745 -267 3779 -233
rect 3813 -267 3847 -233
rect 3881 -267 3915 -233
rect 3949 -267 3983 -233
rect 4017 -267 4051 -233
rect 4085 -267 4119 -233
rect 4153 -267 4187 -233
rect 4221 -267 4255 -233
rect 4289 -267 4323 -233
rect 4357 -267 4391 -233
rect 4425 -267 4459 -233
rect 4493 -267 4527 -233
rect 4561 -267 4595 -233
rect 4629 -267 4663 -233
rect 4697 -267 4731 -233
rect 4765 -267 4799 -233
rect 4833 -267 4867 -233
rect 4901 -267 4935 -233
rect 4969 -267 5003 -233
rect 5037 -267 5071 -233
rect 5105 -267 5139 -233
rect 5173 -267 5207 -233
rect 5241 -267 5275 -233
rect 5309 -267 5343 -233
rect 5377 -267 5411 -233
rect 5445 -267 5479 -233
rect 5513 -267 5547 -233
rect 5581 -267 5615 -233
rect 5649 -267 5683 -233
rect 5717 -267 5751 -233
rect 5785 -267 5819 -233
rect 5853 -267 5887 -233
rect 5921 -267 5955 -233
rect 5989 -267 6023 -233
rect 6057 -267 6091 -233
rect 6125 -267 6159 -233
rect 6193 -267 6227 -233
rect 6261 -267 6295 -233
rect 6329 -267 6363 -233
rect 6397 -267 6431 -233
rect 6465 -267 6499 -233
rect 6533 -267 6567 -233
rect 6601 -267 6635 -233
rect 6669 -267 6703 -233
rect 6737 -267 6771 -233
rect 6805 -267 6839 -233
rect 6873 -267 6907 -233
rect 6941 -267 6975 -233
rect 7009 -267 7043 -233
rect 7077 -267 7111 -233
rect 7145 -267 7179 -233
rect 7213 -267 7247 -233
rect 7281 -267 7315 -233
rect 7349 -267 7383 -233
rect 7417 -267 7451 -233
rect 7485 -267 7519 -233
rect 7553 -267 7587 -233
rect 7621 -267 7655 -233
rect 7689 -267 7723 -233
rect 7757 -267 7791 -233
rect 7825 -267 7859 -233
rect 7893 -267 7927 -233
rect 7961 -267 8000 -233
rect 408 -272 8000 -267
<< psubdiffcont >>
rect 447 -267 481 -233
rect 515 -267 549 -233
rect 583 -267 617 -233
rect 651 -267 685 -233
rect 719 -267 753 -233
rect 787 -267 821 -233
rect 855 -267 889 -233
rect 923 -267 957 -233
rect 991 -267 1025 -233
rect 1059 -267 1093 -233
rect 1127 -267 1161 -233
rect 1195 -267 1229 -233
rect 1263 -267 1297 -233
rect 1331 -267 1365 -233
rect 1399 -267 1433 -233
rect 1467 -267 1501 -233
rect 1535 -267 1569 -233
rect 1603 -267 1637 -233
rect 1671 -267 1705 -233
rect 1739 -267 1773 -233
rect 1807 -267 1841 -233
rect 1875 -267 1909 -233
rect 1943 -267 1977 -233
rect 2011 -267 2045 -233
rect 2079 -267 2113 -233
rect 2147 -267 2181 -233
rect 2215 -267 2249 -233
rect 2283 -267 2317 -233
rect 2351 -267 2385 -233
rect 2419 -267 2453 -233
rect 2487 -267 2521 -233
rect 2555 -267 2589 -233
rect 2623 -267 2657 -233
rect 2691 -267 2725 -233
rect 2759 -267 2793 -233
rect 2827 -267 2861 -233
rect 2895 -267 2929 -233
rect 2963 -267 2997 -233
rect 3031 -267 3065 -233
rect 3099 -267 3133 -233
rect 3167 -267 3201 -233
rect 3235 -267 3269 -233
rect 3303 -267 3337 -233
rect 3371 -267 3405 -233
rect 3439 -267 3473 -233
rect 3507 -267 3541 -233
rect 3575 -267 3609 -233
rect 3643 -267 3677 -233
rect 3711 -267 3745 -233
rect 3779 -267 3813 -233
rect 3847 -267 3881 -233
rect 3915 -267 3949 -233
rect 3983 -267 4017 -233
rect 4051 -267 4085 -233
rect 4119 -267 4153 -233
rect 4187 -267 4221 -233
rect 4255 -267 4289 -233
rect 4323 -267 4357 -233
rect 4391 -267 4425 -233
rect 4459 -267 4493 -233
rect 4527 -267 4561 -233
rect 4595 -267 4629 -233
rect 4663 -267 4697 -233
rect 4731 -267 4765 -233
rect 4799 -267 4833 -233
rect 4867 -267 4901 -233
rect 4935 -267 4969 -233
rect 5003 -267 5037 -233
rect 5071 -267 5105 -233
rect 5139 -267 5173 -233
rect 5207 -267 5241 -233
rect 5275 -267 5309 -233
rect 5343 -267 5377 -233
rect 5411 -267 5445 -233
rect 5479 -267 5513 -233
rect 5547 -267 5581 -233
rect 5615 -267 5649 -233
rect 5683 -267 5717 -233
rect 5751 -267 5785 -233
rect 5819 -267 5853 -233
rect 5887 -267 5921 -233
rect 5955 -267 5989 -233
rect 6023 -267 6057 -233
rect 6091 -267 6125 -233
rect 6159 -267 6193 -233
rect 6227 -267 6261 -233
rect 6295 -267 6329 -233
rect 6363 -267 6397 -233
rect 6431 -267 6465 -233
rect 6499 -267 6533 -233
rect 6567 -267 6601 -233
rect 6635 -267 6669 -233
rect 6703 -267 6737 -233
rect 6771 -267 6805 -233
rect 6839 -267 6873 -233
rect 6907 -267 6941 -233
rect 6975 -267 7009 -233
rect 7043 -267 7077 -233
rect 7111 -267 7145 -233
rect 7179 -267 7213 -233
rect 7247 -267 7281 -233
rect 7315 -267 7349 -233
rect 7383 -267 7417 -233
rect 7451 -267 7485 -233
rect 7519 -267 7553 -233
rect 7587 -267 7621 -233
rect 7655 -267 7689 -233
rect 7723 -267 7757 -233
rect 7791 -267 7825 -233
rect 7859 -267 7893 -233
rect 7927 -267 7961 -233
<< xpolycontact >>
rect 208 1681 278 2113
rect 208 -127 278 305
rect 530 1681 600 2113
rect 530 -127 600 305
rect 852 1681 922 2113
rect 852 -127 922 305
rect 1174 1681 1244 2113
rect 1174 -127 1244 305
rect 1496 1681 1566 2113
rect 1496 -127 1566 305
rect 1818 1681 1888 2113
rect 1818 -127 1888 305
rect 2140 1681 2210 2113
rect 2140 -127 2210 305
rect 2462 1681 2532 2113
rect 2462 -127 2532 305
rect 2784 1681 2854 2113
rect 2784 -127 2854 305
rect 3106 1681 3176 2113
rect 3106 -127 3176 305
rect 3428 1681 3498 2113
rect 3428 -127 3498 305
rect 3750 1681 3820 2113
rect 3750 -127 3820 305
rect 4072 1681 4142 2113
rect 4072 -127 4142 305
rect 4394 1681 4464 2113
rect 4394 -127 4464 305
rect 4716 1681 4786 2113
rect 4716 -127 4786 305
rect 5038 1681 5108 2113
rect 5038 -127 5108 305
rect 5360 1681 5430 2113
rect 5360 -127 5430 305
rect 5682 1681 5752 2113
rect 5682 -127 5752 305
rect 6004 1681 6074 2113
rect 6004 -127 6074 305
rect 6326 1681 6396 2113
rect 6326 -127 6396 305
rect 6648 1681 6718 2113
rect 6648 -127 6718 305
rect 6970 1681 7040 2113
rect 6970 -127 7040 305
rect 7292 1681 7362 2113
rect 7292 -127 7362 305
rect 7614 1681 7684 2113
rect 7614 -127 7684 305
rect 7936 1681 8006 2113
rect 7936 -127 8006 305
rect 204 -807 274 -375
rect 204 -2615 274 -2183
rect 526 -807 596 -375
rect 526 -2615 596 -2183
rect 848 -807 918 -375
rect 848 -2615 918 -2183
rect 1170 -807 1240 -375
rect 1170 -2615 1240 -2183
rect 1492 -807 1562 -375
rect 1492 -2615 1562 -2183
rect 1814 -807 1884 -375
rect 1814 -2615 1884 -2183
rect 2136 -807 2206 -375
rect 2136 -2615 2206 -2183
rect 2458 -807 2528 -375
rect 2458 -2615 2528 -2183
rect 2780 -807 2850 -375
rect 2780 -2615 2850 -2183
rect 3102 -807 3172 -375
rect 3102 -2615 3172 -2183
rect 3424 -807 3494 -375
rect 3424 -2615 3494 -2183
rect 3746 -807 3816 -375
rect 3746 -2615 3816 -2183
rect 4068 -807 4138 -375
rect 4068 -2615 4138 -2183
rect 4390 -807 4460 -375
rect 4390 -2615 4460 -2183
rect 4712 -807 4782 -375
rect 4712 -2615 4782 -2183
rect 5034 -807 5104 -375
rect 5034 -2615 5104 -2183
rect 5356 -807 5426 -375
rect 5356 -2615 5426 -2183
rect 5678 -807 5748 -375
rect 5678 -2615 5748 -2183
rect 6000 -807 6070 -375
rect 6000 -2615 6070 -2183
rect 6322 -807 6392 -375
rect 6322 -2615 6392 -2183
rect 6644 -807 6714 -375
rect 6644 -2615 6714 -2183
rect 6966 -807 7036 -375
rect 6966 -2615 7036 -2183
rect 7288 -807 7358 -375
rect 7288 -2615 7358 -2183
rect 7610 -807 7680 -375
rect 7610 -2615 7680 -2183
rect 7932 -807 8002 -375
rect 7932 -2615 8002 -2183
<< xpolyres >>
rect 208 305 278 1681
rect 530 305 600 1681
rect 852 305 922 1681
rect 1174 305 1244 1681
rect 1496 305 1566 1681
rect 1818 305 1888 1681
rect 2140 305 2210 1681
rect 2462 305 2532 1681
rect 2784 305 2854 1681
rect 3106 305 3176 1681
rect 3428 305 3498 1681
rect 3750 305 3820 1681
rect 4072 305 4142 1681
rect 4394 305 4464 1681
rect 4716 305 4786 1681
rect 5038 305 5108 1681
rect 5360 305 5430 1681
rect 5682 305 5752 1681
rect 6004 305 6074 1681
rect 6326 305 6396 1681
rect 6648 305 6718 1681
rect 6970 305 7040 1681
rect 7292 305 7362 1681
rect 7614 305 7684 1681
rect 7936 305 8006 1681
rect 204 -2183 274 -807
rect 526 -2183 596 -807
rect 848 -2183 918 -807
rect 1170 -2183 1240 -807
rect 1492 -2183 1562 -807
rect 1814 -2183 1884 -807
rect 2136 -2183 2206 -807
rect 2458 -2183 2528 -807
rect 2780 -2183 2850 -807
rect 3102 -2183 3172 -807
rect 3424 -2183 3494 -807
rect 3746 -2183 3816 -807
rect 4068 -2183 4138 -807
rect 4390 -2183 4460 -807
rect 4712 -2183 4782 -807
rect 5034 -2183 5104 -807
rect 5356 -2183 5426 -807
rect 5678 -2183 5748 -807
rect 6000 -2183 6070 -807
rect 6322 -2183 6392 -807
rect 6644 -2183 6714 -807
rect 6966 -2183 7036 -807
rect 7288 -2183 7358 -807
rect 7610 -2183 7680 -807
rect 7932 -2183 8002 -807
<< locali >>
rect 416 -233 7992 -228
rect 416 -267 447 -233
rect 481 -267 515 -233
rect 549 -267 583 -233
rect 617 -267 651 -233
rect 685 -267 719 -233
rect 753 -267 787 -233
rect 821 -267 855 -233
rect 889 -267 923 -233
rect 957 -267 991 -233
rect 1025 -267 1059 -233
rect 1093 -267 1127 -233
rect 1161 -267 1195 -233
rect 1229 -267 1263 -233
rect 1297 -267 1331 -233
rect 1365 -267 1399 -233
rect 1433 -267 1467 -233
rect 1501 -267 1535 -233
rect 1569 -267 1603 -233
rect 1637 -267 1671 -233
rect 1705 -267 1739 -233
rect 1773 -267 1807 -233
rect 1841 -267 1875 -233
rect 1909 -267 1943 -233
rect 1977 -267 2011 -233
rect 2045 -267 2079 -233
rect 2113 -267 2147 -233
rect 2181 -267 2215 -233
rect 2249 -267 2283 -233
rect 2317 -267 2351 -233
rect 2385 -267 2419 -233
rect 2453 -267 2487 -233
rect 2521 -267 2555 -233
rect 2589 -267 2623 -233
rect 2657 -267 2691 -233
rect 2725 -267 2759 -233
rect 2793 -267 2827 -233
rect 2861 -267 2895 -233
rect 2929 -267 2963 -233
rect 2997 -267 3031 -233
rect 3065 -267 3099 -233
rect 3133 -267 3167 -233
rect 3201 -267 3235 -233
rect 3269 -267 3303 -233
rect 3337 -267 3371 -233
rect 3405 -267 3439 -233
rect 3473 -267 3507 -233
rect 3541 -267 3575 -233
rect 3609 -267 3643 -233
rect 3677 -267 3711 -233
rect 3745 -267 3779 -233
rect 3813 -267 3847 -233
rect 3881 -267 3915 -233
rect 3949 -267 3983 -233
rect 4017 -267 4051 -233
rect 4085 -267 4119 -233
rect 4153 -267 4187 -233
rect 4221 -267 4255 -233
rect 4289 -267 4323 -233
rect 4357 -267 4391 -233
rect 4425 -267 4459 -233
rect 4493 -267 4527 -233
rect 4561 -267 4595 -233
rect 4629 -267 4663 -233
rect 4697 -267 4731 -233
rect 4765 -267 4799 -233
rect 4833 -267 4867 -233
rect 4901 -267 4935 -233
rect 4969 -267 5003 -233
rect 5037 -267 5071 -233
rect 5105 -267 5139 -233
rect 5173 -267 5207 -233
rect 5241 -267 5275 -233
rect 5309 -267 5343 -233
rect 5377 -267 5411 -233
rect 5445 -267 5479 -233
rect 5513 -267 5547 -233
rect 5581 -267 5615 -233
rect 5649 -267 5683 -233
rect 5717 -267 5751 -233
rect 5785 -267 5819 -233
rect 5853 -267 5887 -233
rect 5921 -267 5955 -233
rect 5989 -267 6023 -233
rect 6057 -267 6091 -233
rect 6125 -267 6159 -233
rect 6193 -267 6227 -233
rect 6261 -267 6295 -233
rect 6329 -267 6363 -233
rect 6397 -267 6431 -233
rect 6465 -267 6499 -233
rect 6533 -267 6567 -233
rect 6601 -267 6635 -233
rect 6669 -267 6703 -233
rect 6737 -267 6771 -233
rect 6805 -267 6839 -233
rect 6873 -267 6907 -233
rect 6941 -267 6975 -233
rect 7009 -267 7043 -233
rect 7077 -267 7111 -233
rect 7145 -267 7179 -233
rect 7213 -267 7247 -233
rect 7281 -267 7315 -233
rect 7349 -267 7383 -233
rect 7417 -267 7451 -233
rect 7485 -267 7519 -233
rect 7553 -267 7587 -233
rect 7621 -267 7655 -233
rect 7689 -267 7723 -233
rect 7757 -267 7791 -233
rect 7825 -267 7859 -233
rect 7893 -267 7927 -233
rect 7961 -267 7992 -233
rect 416 -272 7992 -267
<< viali >>
rect 226 2059 260 2093
rect 226 1987 260 2021
rect 226 1915 260 1949
rect 226 1843 260 1877
rect 226 1771 260 1805
rect 226 1699 260 1733
rect 548 2059 582 2093
rect 548 1987 582 2021
rect 548 1915 582 1949
rect 548 1843 582 1877
rect 548 1771 582 1805
rect 548 1699 582 1733
rect 870 2059 904 2093
rect 870 1987 904 2021
rect 870 1915 904 1949
rect 870 1843 904 1877
rect 870 1771 904 1805
rect 870 1699 904 1733
rect 1192 2059 1226 2093
rect 1192 1987 1226 2021
rect 1192 1915 1226 1949
rect 1192 1843 1226 1877
rect 1192 1771 1226 1805
rect 1192 1699 1226 1733
rect 1514 2059 1548 2093
rect 1514 1987 1548 2021
rect 1514 1915 1548 1949
rect 1514 1843 1548 1877
rect 1514 1771 1548 1805
rect 1514 1699 1548 1733
rect 1836 2059 1870 2093
rect 1836 1987 1870 2021
rect 1836 1915 1870 1949
rect 1836 1843 1870 1877
rect 1836 1771 1870 1805
rect 1836 1699 1870 1733
rect 2158 2059 2192 2093
rect 2158 1987 2192 2021
rect 2158 1915 2192 1949
rect 2158 1843 2192 1877
rect 2158 1771 2192 1805
rect 2158 1699 2192 1733
rect 2480 2059 2514 2093
rect 2480 1987 2514 2021
rect 2480 1915 2514 1949
rect 2480 1843 2514 1877
rect 2480 1771 2514 1805
rect 2480 1699 2514 1733
rect 2802 2059 2836 2093
rect 2802 1987 2836 2021
rect 2802 1915 2836 1949
rect 2802 1843 2836 1877
rect 2802 1771 2836 1805
rect 2802 1699 2836 1733
rect 3124 2059 3158 2093
rect 3124 1987 3158 2021
rect 3124 1915 3158 1949
rect 3124 1843 3158 1877
rect 3124 1771 3158 1805
rect 3124 1699 3158 1733
rect 3446 2059 3480 2093
rect 3446 1987 3480 2021
rect 3446 1915 3480 1949
rect 3446 1843 3480 1877
rect 3446 1771 3480 1805
rect 3446 1699 3480 1733
rect 3768 2059 3802 2093
rect 3768 1987 3802 2021
rect 3768 1915 3802 1949
rect 3768 1843 3802 1877
rect 3768 1771 3802 1805
rect 3768 1699 3802 1733
rect 4090 2059 4124 2093
rect 4090 1987 4124 2021
rect 4090 1915 4124 1949
rect 4090 1843 4124 1877
rect 4090 1771 4124 1805
rect 4090 1699 4124 1733
rect 4412 2059 4446 2093
rect 4412 1987 4446 2021
rect 4412 1915 4446 1949
rect 4412 1843 4446 1877
rect 4412 1771 4446 1805
rect 4412 1699 4446 1733
rect 4734 2059 4768 2093
rect 4734 1987 4768 2021
rect 4734 1915 4768 1949
rect 4734 1843 4768 1877
rect 4734 1771 4768 1805
rect 4734 1699 4768 1733
rect 5056 2059 5090 2093
rect 5056 1987 5090 2021
rect 5056 1915 5090 1949
rect 5056 1843 5090 1877
rect 5056 1771 5090 1805
rect 5056 1699 5090 1733
rect 5378 2059 5412 2093
rect 5378 1987 5412 2021
rect 5378 1915 5412 1949
rect 5378 1843 5412 1877
rect 5378 1771 5412 1805
rect 5378 1699 5412 1733
rect 5700 2059 5734 2093
rect 5700 1987 5734 2021
rect 5700 1915 5734 1949
rect 5700 1843 5734 1877
rect 5700 1771 5734 1805
rect 5700 1699 5734 1733
rect 6022 2059 6056 2093
rect 6022 1987 6056 2021
rect 6022 1915 6056 1949
rect 6022 1843 6056 1877
rect 6022 1771 6056 1805
rect 6022 1699 6056 1733
rect 6344 2059 6378 2093
rect 6344 1987 6378 2021
rect 6344 1915 6378 1949
rect 6344 1843 6378 1877
rect 6344 1771 6378 1805
rect 6344 1699 6378 1733
rect 6666 2059 6700 2093
rect 6666 1987 6700 2021
rect 6666 1915 6700 1949
rect 6666 1843 6700 1877
rect 6666 1771 6700 1805
rect 6666 1699 6700 1733
rect 6988 2059 7022 2093
rect 6988 1987 7022 2021
rect 6988 1915 7022 1949
rect 6988 1843 7022 1877
rect 6988 1771 7022 1805
rect 6988 1699 7022 1733
rect 7310 2059 7344 2093
rect 7310 1987 7344 2021
rect 7310 1915 7344 1949
rect 7310 1843 7344 1877
rect 7310 1771 7344 1805
rect 7310 1699 7344 1733
rect 7632 2059 7666 2093
rect 7632 1987 7666 2021
rect 7632 1915 7666 1949
rect 7632 1843 7666 1877
rect 7632 1771 7666 1805
rect 7632 1699 7666 1733
rect 7954 2059 7988 2093
rect 7954 1987 7988 2021
rect 7954 1915 7988 1949
rect 7954 1843 7988 1877
rect 7954 1771 7988 1805
rect 7954 1699 7988 1733
rect 226 252 260 286
rect 226 180 260 214
rect 226 108 260 142
rect 226 36 260 70
rect 226 -36 260 -2
rect 226 -108 260 -74
rect 548 252 582 286
rect 548 180 582 214
rect 548 108 582 142
rect 548 36 582 70
rect 548 -36 582 -2
rect 548 -108 582 -74
rect 870 252 904 286
rect 870 180 904 214
rect 870 108 904 142
rect 870 36 904 70
rect 870 -36 904 -2
rect 870 -108 904 -74
rect 1192 252 1226 286
rect 1192 180 1226 214
rect 1192 108 1226 142
rect 1192 36 1226 70
rect 1192 -36 1226 -2
rect 1192 -108 1226 -74
rect 1514 252 1548 286
rect 1514 180 1548 214
rect 1514 108 1548 142
rect 1514 36 1548 70
rect 1514 -36 1548 -2
rect 1514 -108 1548 -74
rect 1836 252 1870 286
rect 1836 180 1870 214
rect 1836 108 1870 142
rect 1836 36 1870 70
rect 1836 -36 1870 -2
rect 1836 -108 1870 -74
rect 2158 252 2192 286
rect 2158 180 2192 214
rect 2158 108 2192 142
rect 2158 36 2192 70
rect 2158 -36 2192 -2
rect 2158 -108 2192 -74
rect 2480 252 2514 286
rect 2480 180 2514 214
rect 2480 108 2514 142
rect 2480 36 2514 70
rect 2480 -36 2514 -2
rect 2480 -108 2514 -74
rect 2802 252 2836 286
rect 2802 180 2836 214
rect 2802 108 2836 142
rect 2802 36 2836 70
rect 2802 -36 2836 -2
rect 2802 -108 2836 -74
rect 3124 252 3158 286
rect 3124 180 3158 214
rect 3124 108 3158 142
rect 3124 36 3158 70
rect 3124 -36 3158 -2
rect 3124 -108 3158 -74
rect 3446 252 3480 286
rect 3446 180 3480 214
rect 3446 108 3480 142
rect 3446 36 3480 70
rect 3446 -36 3480 -2
rect 3446 -108 3480 -74
rect 3768 252 3802 286
rect 3768 180 3802 214
rect 3768 108 3802 142
rect 3768 36 3802 70
rect 3768 -36 3802 -2
rect 3768 -108 3802 -74
rect 4090 252 4124 286
rect 4090 180 4124 214
rect 4090 108 4124 142
rect 4090 36 4124 70
rect 4090 -36 4124 -2
rect 4090 -108 4124 -74
rect 4412 252 4446 286
rect 4412 180 4446 214
rect 4412 108 4446 142
rect 4412 36 4446 70
rect 4412 -36 4446 -2
rect 4412 -108 4446 -74
rect 4734 252 4768 286
rect 4734 180 4768 214
rect 4734 108 4768 142
rect 4734 36 4768 70
rect 4734 -36 4768 -2
rect 4734 -108 4768 -74
rect 5056 252 5090 286
rect 5056 180 5090 214
rect 5056 108 5090 142
rect 5056 36 5090 70
rect 5056 -36 5090 -2
rect 5056 -108 5090 -74
rect 5378 252 5412 286
rect 5378 180 5412 214
rect 5378 108 5412 142
rect 5378 36 5412 70
rect 5378 -36 5412 -2
rect 5378 -108 5412 -74
rect 5700 252 5734 286
rect 5700 180 5734 214
rect 5700 108 5734 142
rect 5700 36 5734 70
rect 5700 -36 5734 -2
rect 5700 -108 5734 -74
rect 6022 252 6056 286
rect 6022 180 6056 214
rect 6022 108 6056 142
rect 6022 36 6056 70
rect 6022 -36 6056 -2
rect 6022 -108 6056 -74
rect 6344 252 6378 286
rect 6344 180 6378 214
rect 6344 108 6378 142
rect 6344 36 6378 70
rect 6344 -36 6378 -2
rect 6344 -108 6378 -74
rect 6666 252 6700 286
rect 6666 180 6700 214
rect 6666 108 6700 142
rect 6666 36 6700 70
rect 6666 -36 6700 -2
rect 6666 -108 6700 -74
rect 6988 252 7022 286
rect 6988 180 7022 214
rect 6988 108 7022 142
rect 6988 36 7022 70
rect 6988 -36 7022 -2
rect 6988 -108 7022 -74
rect 7310 252 7344 286
rect 7310 180 7344 214
rect 7310 108 7344 142
rect 7310 36 7344 70
rect 7310 -36 7344 -2
rect 7310 -108 7344 -74
rect 7632 252 7666 286
rect 7632 180 7666 214
rect 7632 108 7666 142
rect 7632 36 7666 70
rect 7632 -36 7666 -2
rect 7632 -108 7666 -74
rect 7954 252 7988 286
rect 7954 180 7988 214
rect 7954 108 7988 142
rect 7954 36 7988 70
rect 7954 -36 7988 -2
rect 7954 -108 7988 -74
rect 222 -429 256 -395
rect 222 -501 256 -467
rect 222 -573 256 -539
rect 222 -645 256 -611
rect 222 -717 256 -683
rect 222 -789 256 -755
rect 544 -429 578 -395
rect 544 -501 578 -467
rect 544 -573 578 -539
rect 544 -645 578 -611
rect 544 -717 578 -683
rect 544 -789 578 -755
rect 866 -429 900 -395
rect 866 -501 900 -467
rect 866 -573 900 -539
rect 866 -645 900 -611
rect 866 -717 900 -683
rect 866 -789 900 -755
rect 1188 -429 1222 -395
rect 1188 -501 1222 -467
rect 1188 -573 1222 -539
rect 1188 -645 1222 -611
rect 1188 -717 1222 -683
rect 1188 -789 1222 -755
rect 1510 -429 1544 -395
rect 1510 -501 1544 -467
rect 1510 -573 1544 -539
rect 1510 -645 1544 -611
rect 1510 -717 1544 -683
rect 1510 -789 1544 -755
rect 1832 -429 1866 -395
rect 1832 -501 1866 -467
rect 1832 -573 1866 -539
rect 1832 -645 1866 -611
rect 1832 -717 1866 -683
rect 1832 -789 1866 -755
rect 2154 -429 2188 -395
rect 2154 -501 2188 -467
rect 2154 -573 2188 -539
rect 2154 -645 2188 -611
rect 2154 -717 2188 -683
rect 2154 -789 2188 -755
rect 2476 -429 2510 -395
rect 2476 -501 2510 -467
rect 2476 -573 2510 -539
rect 2476 -645 2510 -611
rect 2476 -717 2510 -683
rect 2476 -789 2510 -755
rect 2798 -429 2832 -395
rect 2798 -501 2832 -467
rect 2798 -573 2832 -539
rect 2798 -645 2832 -611
rect 2798 -717 2832 -683
rect 2798 -789 2832 -755
rect 3120 -429 3154 -395
rect 3120 -501 3154 -467
rect 3120 -573 3154 -539
rect 3120 -645 3154 -611
rect 3120 -717 3154 -683
rect 3120 -789 3154 -755
rect 3442 -429 3476 -395
rect 3442 -501 3476 -467
rect 3442 -573 3476 -539
rect 3442 -645 3476 -611
rect 3442 -717 3476 -683
rect 3442 -789 3476 -755
rect 3764 -429 3798 -395
rect 3764 -501 3798 -467
rect 3764 -573 3798 -539
rect 3764 -645 3798 -611
rect 3764 -717 3798 -683
rect 3764 -789 3798 -755
rect 4086 -429 4120 -395
rect 4086 -501 4120 -467
rect 4086 -573 4120 -539
rect 4086 -645 4120 -611
rect 4086 -717 4120 -683
rect 4086 -789 4120 -755
rect 4408 -429 4442 -395
rect 4408 -501 4442 -467
rect 4408 -573 4442 -539
rect 4408 -645 4442 -611
rect 4408 -717 4442 -683
rect 4408 -789 4442 -755
rect 4730 -429 4764 -395
rect 4730 -501 4764 -467
rect 4730 -573 4764 -539
rect 4730 -645 4764 -611
rect 4730 -717 4764 -683
rect 4730 -789 4764 -755
rect 5052 -429 5086 -395
rect 5052 -501 5086 -467
rect 5052 -573 5086 -539
rect 5052 -645 5086 -611
rect 5052 -717 5086 -683
rect 5052 -789 5086 -755
rect 5374 -429 5408 -395
rect 5374 -501 5408 -467
rect 5374 -573 5408 -539
rect 5374 -645 5408 -611
rect 5374 -717 5408 -683
rect 5374 -789 5408 -755
rect 5696 -429 5730 -395
rect 5696 -501 5730 -467
rect 5696 -573 5730 -539
rect 5696 -645 5730 -611
rect 5696 -717 5730 -683
rect 5696 -789 5730 -755
rect 6018 -429 6052 -395
rect 6018 -501 6052 -467
rect 6018 -573 6052 -539
rect 6018 -645 6052 -611
rect 6018 -717 6052 -683
rect 6018 -789 6052 -755
rect 6340 -429 6374 -395
rect 6340 -501 6374 -467
rect 6340 -573 6374 -539
rect 6340 -645 6374 -611
rect 6340 -717 6374 -683
rect 6340 -789 6374 -755
rect 6662 -429 6696 -395
rect 6662 -501 6696 -467
rect 6662 -573 6696 -539
rect 6662 -645 6696 -611
rect 6662 -717 6696 -683
rect 6662 -789 6696 -755
rect 6984 -429 7018 -395
rect 6984 -501 7018 -467
rect 6984 -573 7018 -539
rect 6984 -645 7018 -611
rect 6984 -717 7018 -683
rect 6984 -789 7018 -755
rect 7306 -429 7340 -395
rect 7306 -501 7340 -467
rect 7306 -573 7340 -539
rect 7306 -645 7340 -611
rect 7306 -717 7340 -683
rect 7306 -789 7340 -755
rect 7628 -429 7662 -395
rect 7628 -501 7662 -467
rect 7628 -573 7662 -539
rect 7628 -645 7662 -611
rect 7628 -717 7662 -683
rect 7628 -789 7662 -755
rect 7950 -429 7984 -395
rect 7950 -501 7984 -467
rect 7950 -573 7984 -539
rect 7950 -645 7984 -611
rect 7950 -717 7984 -683
rect 7950 -789 7984 -755
rect 222 -2236 256 -2202
rect 222 -2308 256 -2274
rect 222 -2380 256 -2346
rect 222 -2452 256 -2418
rect 222 -2524 256 -2490
rect 222 -2596 256 -2562
rect 544 -2236 578 -2202
rect 544 -2308 578 -2274
rect 544 -2380 578 -2346
rect 544 -2452 578 -2418
rect 544 -2524 578 -2490
rect 544 -2596 578 -2562
rect 866 -2236 900 -2202
rect 866 -2308 900 -2274
rect 866 -2380 900 -2346
rect 866 -2452 900 -2418
rect 866 -2524 900 -2490
rect 866 -2596 900 -2562
rect 1188 -2236 1222 -2202
rect 1188 -2308 1222 -2274
rect 1188 -2380 1222 -2346
rect 1188 -2452 1222 -2418
rect 1188 -2524 1222 -2490
rect 1188 -2596 1222 -2562
rect 1510 -2236 1544 -2202
rect 1510 -2308 1544 -2274
rect 1510 -2380 1544 -2346
rect 1510 -2452 1544 -2418
rect 1510 -2524 1544 -2490
rect 1510 -2596 1544 -2562
rect 1832 -2236 1866 -2202
rect 1832 -2308 1866 -2274
rect 1832 -2380 1866 -2346
rect 1832 -2452 1866 -2418
rect 1832 -2524 1866 -2490
rect 1832 -2596 1866 -2562
rect 2154 -2236 2188 -2202
rect 2154 -2308 2188 -2274
rect 2154 -2380 2188 -2346
rect 2154 -2452 2188 -2418
rect 2154 -2524 2188 -2490
rect 2154 -2596 2188 -2562
rect 2476 -2236 2510 -2202
rect 2476 -2308 2510 -2274
rect 2476 -2380 2510 -2346
rect 2476 -2452 2510 -2418
rect 2476 -2524 2510 -2490
rect 2476 -2596 2510 -2562
rect 2798 -2236 2832 -2202
rect 2798 -2308 2832 -2274
rect 2798 -2380 2832 -2346
rect 2798 -2452 2832 -2418
rect 2798 -2524 2832 -2490
rect 2798 -2596 2832 -2562
rect 3120 -2236 3154 -2202
rect 3120 -2308 3154 -2274
rect 3120 -2380 3154 -2346
rect 3120 -2452 3154 -2418
rect 3120 -2524 3154 -2490
rect 3120 -2596 3154 -2562
rect 3442 -2236 3476 -2202
rect 3442 -2308 3476 -2274
rect 3442 -2380 3476 -2346
rect 3442 -2452 3476 -2418
rect 3442 -2524 3476 -2490
rect 3442 -2596 3476 -2562
rect 3764 -2236 3798 -2202
rect 3764 -2308 3798 -2274
rect 3764 -2380 3798 -2346
rect 3764 -2452 3798 -2418
rect 3764 -2524 3798 -2490
rect 3764 -2596 3798 -2562
rect 4086 -2236 4120 -2202
rect 4086 -2308 4120 -2274
rect 4086 -2380 4120 -2346
rect 4086 -2452 4120 -2418
rect 4086 -2524 4120 -2490
rect 4086 -2596 4120 -2562
rect 4408 -2236 4442 -2202
rect 4408 -2308 4442 -2274
rect 4408 -2380 4442 -2346
rect 4408 -2452 4442 -2418
rect 4408 -2524 4442 -2490
rect 4408 -2596 4442 -2562
rect 4730 -2236 4764 -2202
rect 4730 -2308 4764 -2274
rect 4730 -2380 4764 -2346
rect 4730 -2452 4764 -2418
rect 4730 -2524 4764 -2490
rect 4730 -2596 4764 -2562
rect 5052 -2236 5086 -2202
rect 5052 -2308 5086 -2274
rect 5052 -2380 5086 -2346
rect 5052 -2452 5086 -2418
rect 5052 -2524 5086 -2490
rect 5052 -2596 5086 -2562
rect 5374 -2236 5408 -2202
rect 5374 -2308 5408 -2274
rect 5374 -2380 5408 -2346
rect 5374 -2452 5408 -2418
rect 5374 -2524 5408 -2490
rect 5374 -2596 5408 -2562
rect 5696 -2236 5730 -2202
rect 5696 -2308 5730 -2274
rect 5696 -2380 5730 -2346
rect 5696 -2452 5730 -2418
rect 5696 -2524 5730 -2490
rect 5696 -2596 5730 -2562
rect 6018 -2236 6052 -2202
rect 6018 -2308 6052 -2274
rect 6018 -2380 6052 -2346
rect 6018 -2452 6052 -2418
rect 6018 -2524 6052 -2490
rect 6018 -2596 6052 -2562
rect 6340 -2236 6374 -2202
rect 6340 -2308 6374 -2274
rect 6340 -2380 6374 -2346
rect 6340 -2452 6374 -2418
rect 6340 -2524 6374 -2490
rect 6340 -2596 6374 -2562
rect 6662 -2236 6696 -2202
rect 6662 -2308 6696 -2274
rect 6662 -2380 6696 -2346
rect 6662 -2452 6696 -2418
rect 6662 -2524 6696 -2490
rect 6662 -2596 6696 -2562
rect 6984 -2236 7018 -2202
rect 6984 -2308 7018 -2274
rect 6984 -2380 7018 -2346
rect 6984 -2452 7018 -2418
rect 6984 -2524 7018 -2490
rect 6984 -2596 7018 -2562
rect 7306 -2236 7340 -2202
rect 7306 -2308 7340 -2274
rect 7306 -2380 7340 -2346
rect 7306 -2452 7340 -2418
rect 7306 -2524 7340 -2490
rect 7306 -2596 7340 -2562
rect 7628 -2236 7662 -2202
rect 7628 -2308 7662 -2274
rect 7628 -2380 7662 -2346
rect 7628 -2452 7662 -2418
rect 7628 -2524 7662 -2490
rect 7628 -2596 7662 -2562
rect 7950 -2236 7984 -2202
rect 7950 -2308 7984 -2274
rect 7950 -2380 7984 -2346
rect 7950 -2452 7984 -2418
rect 7950 -2524 7984 -2490
rect 7950 -2596 7984 -2562
<< metal1 >>
rect 7212 2509 8012 2542
rect 7212 2329 7267 2509
rect 7959 2329 8012 2509
rect 7212 2302 8012 2329
rect 208 2093 600 2114
rect 208 2059 226 2093
rect 260 2059 548 2093
rect 582 2059 600 2093
rect 208 2021 600 2059
rect 208 1987 226 2021
rect 260 1987 548 2021
rect 582 1987 600 2021
rect 208 1949 600 1987
rect 208 1915 226 1949
rect 260 1915 548 1949
rect 582 1915 600 1949
rect 208 1877 600 1915
rect 208 1843 226 1877
rect 260 1843 548 1877
rect 582 1843 600 1877
rect 208 1805 600 1843
rect 208 1771 226 1805
rect 260 1771 548 1805
rect 582 1771 600 1805
rect 208 1733 600 1771
rect 208 1699 226 1733
rect 260 1699 548 1733
rect 582 1699 600 1733
rect 208 1680 600 1699
rect 852 2093 1244 2114
rect 852 2059 870 2093
rect 904 2059 1192 2093
rect 1226 2059 1244 2093
rect 852 2021 1244 2059
rect 852 1987 870 2021
rect 904 1987 1192 2021
rect 1226 1987 1244 2021
rect 852 1949 1244 1987
rect 852 1915 870 1949
rect 904 1915 1192 1949
rect 1226 1915 1244 1949
rect 852 1877 1244 1915
rect 852 1843 870 1877
rect 904 1843 1192 1877
rect 1226 1843 1244 1877
rect 852 1805 1244 1843
rect 852 1771 870 1805
rect 904 1771 1192 1805
rect 1226 1771 1244 1805
rect 852 1733 1244 1771
rect 852 1699 870 1733
rect 904 1699 1192 1733
rect 1226 1699 1244 1733
rect 852 1680 1244 1699
rect 1496 2093 1888 2114
rect 1496 2059 1514 2093
rect 1548 2059 1836 2093
rect 1870 2059 1888 2093
rect 1496 2021 1888 2059
rect 1496 1987 1514 2021
rect 1548 1987 1836 2021
rect 1870 1987 1888 2021
rect 1496 1949 1888 1987
rect 1496 1915 1514 1949
rect 1548 1915 1836 1949
rect 1870 1915 1888 1949
rect 1496 1877 1888 1915
rect 1496 1843 1514 1877
rect 1548 1843 1836 1877
rect 1870 1843 1888 1877
rect 1496 1805 1888 1843
rect 1496 1771 1514 1805
rect 1548 1771 1836 1805
rect 1870 1771 1888 1805
rect 1496 1733 1888 1771
rect 1496 1699 1514 1733
rect 1548 1699 1836 1733
rect 1870 1699 1888 1733
rect 1496 1680 1888 1699
rect 2140 2093 2532 2114
rect 2140 2059 2158 2093
rect 2192 2059 2480 2093
rect 2514 2059 2532 2093
rect 2140 2021 2532 2059
rect 2140 1987 2158 2021
rect 2192 1987 2480 2021
rect 2514 1987 2532 2021
rect 2140 1949 2532 1987
rect 2140 1915 2158 1949
rect 2192 1915 2480 1949
rect 2514 1915 2532 1949
rect 2140 1877 2532 1915
rect 2140 1843 2158 1877
rect 2192 1843 2480 1877
rect 2514 1843 2532 1877
rect 2140 1805 2532 1843
rect 2140 1771 2158 1805
rect 2192 1771 2480 1805
rect 2514 1771 2532 1805
rect 2140 1733 2532 1771
rect 2140 1699 2158 1733
rect 2192 1699 2480 1733
rect 2514 1699 2532 1733
rect 2140 1680 2532 1699
rect 2784 2093 3176 2114
rect 2784 2059 2802 2093
rect 2836 2059 3124 2093
rect 3158 2059 3176 2093
rect 2784 2021 3176 2059
rect 2784 1987 2802 2021
rect 2836 1987 3124 2021
rect 3158 1987 3176 2021
rect 2784 1949 3176 1987
rect 2784 1915 2802 1949
rect 2836 1915 3124 1949
rect 3158 1915 3176 1949
rect 2784 1877 3176 1915
rect 2784 1843 2802 1877
rect 2836 1843 3124 1877
rect 3158 1843 3176 1877
rect 2784 1805 3176 1843
rect 2784 1771 2802 1805
rect 2836 1771 3124 1805
rect 3158 1771 3176 1805
rect 2784 1733 3176 1771
rect 2784 1699 2802 1733
rect 2836 1699 3124 1733
rect 3158 1699 3176 1733
rect 2784 1680 3176 1699
rect 3428 2093 3820 2114
rect 3428 2059 3446 2093
rect 3480 2059 3768 2093
rect 3802 2059 3820 2093
rect 3428 2021 3820 2059
rect 3428 1987 3446 2021
rect 3480 1987 3768 2021
rect 3802 1987 3820 2021
rect 3428 1949 3820 1987
rect 3428 1915 3446 1949
rect 3480 1915 3768 1949
rect 3802 1915 3820 1949
rect 3428 1877 3820 1915
rect 3428 1843 3446 1877
rect 3480 1843 3768 1877
rect 3802 1843 3820 1877
rect 3428 1805 3820 1843
rect 3428 1771 3446 1805
rect 3480 1771 3768 1805
rect 3802 1771 3820 1805
rect 3428 1733 3820 1771
rect 3428 1699 3446 1733
rect 3480 1699 3768 1733
rect 3802 1699 3820 1733
rect 3428 1680 3820 1699
rect 4072 2093 4464 2114
rect 4072 2059 4090 2093
rect 4124 2059 4412 2093
rect 4446 2059 4464 2093
rect 4072 2021 4464 2059
rect 4072 1987 4090 2021
rect 4124 1987 4412 2021
rect 4446 1987 4464 2021
rect 4072 1949 4464 1987
rect 4072 1915 4090 1949
rect 4124 1915 4412 1949
rect 4446 1915 4464 1949
rect 4072 1877 4464 1915
rect 4072 1843 4090 1877
rect 4124 1843 4412 1877
rect 4446 1843 4464 1877
rect 4072 1805 4464 1843
rect 4072 1771 4090 1805
rect 4124 1771 4412 1805
rect 4446 1771 4464 1805
rect 4072 1733 4464 1771
rect 4072 1699 4090 1733
rect 4124 1699 4412 1733
rect 4446 1699 4464 1733
rect 4072 1680 4464 1699
rect 4716 2093 5108 2114
rect 4716 2059 4734 2093
rect 4768 2059 5056 2093
rect 5090 2059 5108 2093
rect 4716 2021 5108 2059
rect 4716 1987 4734 2021
rect 4768 1987 5056 2021
rect 5090 1987 5108 2021
rect 4716 1949 5108 1987
rect 4716 1915 4734 1949
rect 4768 1915 5056 1949
rect 5090 1915 5108 1949
rect 4716 1877 5108 1915
rect 4716 1843 4734 1877
rect 4768 1843 5056 1877
rect 5090 1843 5108 1877
rect 4716 1805 5108 1843
rect 4716 1771 4734 1805
rect 4768 1771 5056 1805
rect 5090 1771 5108 1805
rect 4716 1733 5108 1771
rect 4716 1699 4734 1733
rect 4768 1699 5056 1733
rect 5090 1699 5108 1733
rect 4716 1680 5108 1699
rect 5360 2093 5752 2114
rect 5360 2059 5378 2093
rect 5412 2059 5700 2093
rect 5734 2059 5752 2093
rect 5360 2021 5752 2059
rect 5360 1987 5378 2021
rect 5412 1987 5700 2021
rect 5734 1987 5752 2021
rect 5360 1949 5752 1987
rect 5360 1915 5378 1949
rect 5412 1915 5700 1949
rect 5734 1915 5752 1949
rect 5360 1877 5752 1915
rect 5360 1843 5378 1877
rect 5412 1843 5700 1877
rect 5734 1843 5752 1877
rect 5360 1805 5752 1843
rect 5360 1771 5378 1805
rect 5412 1771 5700 1805
rect 5734 1771 5752 1805
rect 5360 1733 5752 1771
rect 5360 1699 5378 1733
rect 5412 1699 5700 1733
rect 5734 1699 5752 1733
rect 5360 1680 5752 1699
rect 6004 2093 6396 2114
rect 6004 2059 6022 2093
rect 6056 2059 6344 2093
rect 6378 2059 6396 2093
rect 6004 2021 6396 2059
rect 6004 1987 6022 2021
rect 6056 1987 6344 2021
rect 6378 1987 6396 2021
rect 6004 1949 6396 1987
rect 6004 1915 6022 1949
rect 6056 1915 6344 1949
rect 6378 1915 6396 1949
rect 6004 1877 6396 1915
rect 6004 1843 6022 1877
rect 6056 1843 6344 1877
rect 6378 1843 6396 1877
rect 6004 1805 6396 1843
rect 6004 1771 6022 1805
rect 6056 1771 6344 1805
rect 6378 1771 6396 1805
rect 6004 1733 6396 1771
rect 6004 1699 6022 1733
rect 6056 1699 6344 1733
rect 6378 1699 6396 1733
rect 6004 1680 6396 1699
rect 6648 2093 7040 2114
rect 6648 2059 6666 2093
rect 6700 2059 6988 2093
rect 7022 2059 7040 2093
rect 6648 2021 7040 2059
rect 6648 1987 6666 2021
rect 6700 1987 6988 2021
rect 7022 1987 7040 2021
rect 6648 1949 7040 1987
rect 6648 1915 6666 1949
rect 6700 1915 6988 1949
rect 7022 1915 7040 1949
rect 6648 1877 7040 1915
rect 6648 1843 6666 1877
rect 6700 1843 6988 1877
rect 7022 1843 7040 1877
rect 6648 1805 7040 1843
rect 6648 1771 6666 1805
rect 6700 1771 6988 1805
rect 7022 1771 7040 1805
rect 6648 1733 7040 1771
rect 6648 1699 6666 1733
rect 6700 1699 6988 1733
rect 7022 1699 7040 1733
rect 6648 1680 7040 1699
rect 7292 2093 7684 2114
rect 7292 2059 7310 2093
rect 7344 2059 7632 2093
rect 7666 2059 7684 2093
rect 7936 2093 8006 2302
rect 7936 2084 7954 2093
rect 7292 2021 7684 2059
rect 7292 1987 7310 2021
rect 7344 1987 7632 2021
rect 7666 1987 7684 2021
rect 7292 1949 7684 1987
rect 7292 1915 7310 1949
rect 7344 1915 7632 1949
rect 7666 1915 7684 1949
rect 7292 1877 7684 1915
rect 7292 1843 7310 1877
rect 7344 1843 7632 1877
rect 7666 1843 7684 1877
rect 7292 1805 7684 1843
rect 7292 1771 7310 1805
rect 7344 1771 7632 1805
rect 7666 1771 7684 1805
rect 7292 1733 7684 1771
rect 7292 1699 7310 1733
rect 7344 1699 7632 1733
rect 7666 1699 7684 1733
rect 7292 1680 7684 1699
rect 7946 2059 7954 2084
rect 7988 2084 8006 2093
rect 7988 2059 7996 2084
rect 7946 2021 7996 2059
rect 7946 1987 7954 2021
rect 7988 1987 7996 2021
rect 7946 1949 7996 1987
rect 7946 1915 7954 1949
rect 7988 1915 7996 1949
rect 7946 1877 7996 1915
rect 7946 1843 7954 1877
rect 7988 1843 7996 1877
rect 7946 1805 7996 1843
rect 7946 1771 7954 1805
rect 7988 1771 7996 1805
rect 7946 1733 7996 1771
rect 7946 1699 7954 1733
rect 7988 1699 7996 1733
rect 7946 1686 7996 1699
rect 0 286 276 306
rect 0 252 226 286
rect 260 252 276 286
rect 0 214 276 252
rect 0 180 226 214
rect 260 180 276 214
rect 0 142 276 180
rect 0 108 226 142
rect 260 108 276 142
rect 0 70 276 108
rect 0 36 226 70
rect 260 36 276 70
rect 0 -2 276 36
rect 0 -36 226 -2
rect 260 -36 276 -2
rect 0 -74 276 -36
rect 0 -108 226 -74
rect 260 -108 276 -74
rect 0 -395 276 -108
rect 530 286 922 306
rect 530 252 548 286
rect 582 252 870 286
rect 904 252 922 286
rect 530 214 922 252
rect 530 180 548 214
rect 582 180 870 214
rect 904 180 922 214
rect 530 142 922 180
rect 530 108 548 142
rect 582 108 870 142
rect 904 108 922 142
rect 530 70 922 108
rect 530 36 548 70
rect 582 36 870 70
rect 904 36 922 70
rect 530 -2 922 36
rect 530 -36 548 -2
rect 582 -36 870 -2
rect 904 -36 922 -2
rect 530 -74 922 -36
rect 530 -108 548 -74
rect 582 -108 870 -74
rect 904 -108 922 -74
rect 530 -128 922 -108
rect 1174 286 1566 306
rect 1174 252 1192 286
rect 1226 252 1514 286
rect 1548 252 1566 286
rect 1174 214 1566 252
rect 1174 180 1192 214
rect 1226 180 1514 214
rect 1548 180 1566 214
rect 1174 142 1566 180
rect 1174 108 1192 142
rect 1226 108 1514 142
rect 1548 108 1566 142
rect 1174 70 1566 108
rect 1174 36 1192 70
rect 1226 36 1514 70
rect 1548 36 1566 70
rect 1174 -2 1566 36
rect 1174 -36 1192 -2
rect 1226 -36 1514 -2
rect 1548 -36 1566 -2
rect 1174 -74 1566 -36
rect 1174 -108 1192 -74
rect 1226 -108 1514 -74
rect 1548 -108 1566 -74
rect 1174 -128 1566 -108
rect 1818 286 2210 306
rect 1818 252 1836 286
rect 1870 252 2158 286
rect 2192 252 2210 286
rect 1818 214 2210 252
rect 1818 180 1836 214
rect 1870 180 2158 214
rect 2192 180 2210 214
rect 1818 142 2210 180
rect 1818 108 1836 142
rect 1870 108 2158 142
rect 2192 108 2210 142
rect 1818 70 2210 108
rect 1818 36 1836 70
rect 1870 36 2158 70
rect 2192 36 2210 70
rect 1818 -2 2210 36
rect 1818 -36 1836 -2
rect 1870 -36 2158 -2
rect 2192 -36 2210 -2
rect 1818 -74 2210 -36
rect 1818 -108 1836 -74
rect 1870 -108 2158 -74
rect 2192 -108 2210 -74
rect 1818 -128 2210 -108
rect 2462 286 2854 306
rect 2462 252 2480 286
rect 2514 252 2802 286
rect 2836 252 2854 286
rect 2462 214 2854 252
rect 2462 180 2480 214
rect 2514 180 2802 214
rect 2836 180 2854 214
rect 2462 142 2854 180
rect 2462 108 2480 142
rect 2514 108 2802 142
rect 2836 108 2854 142
rect 2462 70 2854 108
rect 2462 36 2480 70
rect 2514 36 2802 70
rect 2836 36 2854 70
rect 2462 -2 2854 36
rect 2462 -36 2480 -2
rect 2514 -36 2802 -2
rect 2836 -36 2854 -2
rect 2462 -74 2854 -36
rect 2462 -108 2480 -74
rect 2514 -108 2802 -74
rect 2836 -108 2854 -74
rect 2462 -128 2854 -108
rect 3106 286 3498 306
rect 3106 252 3124 286
rect 3158 252 3446 286
rect 3480 252 3498 286
rect 3106 214 3498 252
rect 3106 180 3124 214
rect 3158 180 3446 214
rect 3480 180 3498 214
rect 3106 142 3498 180
rect 3106 108 3124 142
rect 3158 108 3446 142
rect 3480 108 3498 142
rect 3106 70 3498 108
rect 3106 36 3124 70
rect 3158 36 3446 70
rect 3480 36 3498 70
rect 3106 -2 3498 36
rect 3106 -36 3124 -2
rect 3158 -36 3446 -2
rect 3480 -36 3498 -2
rect 3106 -74 3498 -36
rect 3106 -108 3124 -74
rect 3158 -108 3446 -74
rect 3480 -108 3498 -74
rect 3106 -128 3498 -108
rect 3750 286 4142 306
rect 3750 252 3768 286
rect 3802 252 4090 286
rect 4124 252 4142 286
rect 3750 214 4142 252
rect 3750 180 3768 214
rect 3802 180 4090 214
rect 4124 180 4142 214
rect 3750 142 4142 180
rect 3750 108 3768 142
rect 3802 108 4090 142
rect 4124 108 4142 142
rect 3750 70 4142 108
rect 3750 36 3768 70
rect 3802 36 4090 70
rect 4124 36 4142 70
rect 3750 -2 4142 36
rect 3750 -36 3768 -2
rect 3802 -36 4090 -2
rect 4124 -36 4142 -2
rect 3750 -74 4142 -36
rect 3750 -108 3768 -74
rect 3802 -108 4090 -74
rect 4124 -108 4142 -74
rect 3750 -128 4142 -108
rect 4394 286 4786 306
rect 4394 252 4412 286
rect 4446 252 4734 286
rect 4768 252 4786 286
rect 4394 214 4786 252
rect 4394 180 4412 214
rect 4446 180 4734 214
rect 4768 180 4786 214
rect 4394 142 4786 180
rect 4394 108 4412 142
rect 4446 108 4734 142
rect 4768 108 4786 142
rect 4394 70 4786 108
rect 4394 36 4412 70
rect 4446 36 4734 70
rect 4768 36 4786 70
rect 4394 -2 4786 36
rect 4394 -36 4412 -2
rect 4446 -36 4734 -2
rect 4768 -36 4786 -2
rect 4394 -74 4786 -36
rect 4394 -108 4412 -74
rect 4446 -108 4734 -74
rect 4768 -108 4786 -74
rect 4394 -128 4786 -108
rect 5038 286 5430 306
rect 5038 252 5056 286
rect 5090 252 5378 286
rect 5412 252 5430 286
rect 5038 214 5430 252
rect 5038 180 5056 214
rect 5090 180 5378 214
rect 5412 180 5430 214
rect 5038 142 5430 180
rect 5038 108 5056 142
rect 5090 108 5378 142
rect 5412 108 5430 142
rect 5038 70 5430 108
rect 5038 36 5056 70
rect 5090 36 5378 70
rect 5412 36 5430 70
rect 5038 -2 5430 36
rect 5038 -36 5056 -2
rect 5090 -36 5378 -2
rect 5412 -36 5430 -2
rect 5038 -74 5430 -36
rect 5038 -108 5056 -74
rect 5090 -108 5378 -74
rect 5412 -108 5430 -74
rect 5038 -128 5430 -108
rect 5682 286 6074 306
rect 5682 252 5700 286
rect 5734 252 6022 286
rect 6056 252 6074 286
rect 5682 214 6074 252
rect 5682 180 5700 214
rect 5734 180 6022 214
rect 6056 180 6074 214
rect 5682 142 6074 180
rect 5682 108 5700 142
rect 5734 108 6022 142
rect 6056 108 6074 142
rect 5682 70 6074 108
rect 5682 36 5700 70
rect 5734 36 6022 70
rect 6056 36 6074 70
rect 5682 -2 6074 36
rect 5682 -36 5700 -2
rect 5734 -36 6022 -2
rect 6056 -36 6074 -2
rect 5682 -74 6074 -36
rect 5682 -108 5700 -74
rect 5734 -108 6022 -74
rect 6056 -108 6074 -74
rect 5682 -128 6074 -108
rect 6326 286 6718 306
rect 6326 252 6344 286
rect 6378 252 6666 286
rect 6700 252 6718 286
rect 6326 214 6718 252
rect 6326 180 6344 214
rect 6378 180 6666 214
rect 6700 180 6718 214
rect 6326 142 6718 180
rect 6326 108 6344 142
rect 6378 108 6666 142
rect 6700 108 6718 142
rect 6326 70 6718 108
rect 6326 36 6344 70
rect 6378 36 6666 70
rect 6700 36 6718 70
rect 6326 -2 6718 36
rect 6326 -36 6344 -2
rect 6378 -36 6666 -2
rect 6700 -36 6718 -2
rect 6326 -74 6718 -36
rect 6326 -108 6344 -74
rect 6378 -108 6666 -74
rect 6700 -108 6718 -74
rect 6326 -128 6718 -108
rect 6970 286 7362 306
rect 6970 252 6988 286
rect 7022 252 7310 286
rect 7344 252 7362 286
rect 6970 214 7362 252
rect 6970 180 6988 214
rect 7022 180 7310 214
rect 7344 180 7362 214
rect 6970 142 7362 180
rect 6970 108 6988 142
rect 7022 108 7310 142
rect 7344 108 7362 142
rect 6970 70 7362 108
rect 6970 36 6988 70
rect 7022 36 7310 70
rect 7344 36 7362 70
rect 6970 -2 7362 36
rect 6970 -36 6988 -2
rect 7022 -36 7310 -2
rect 7344 -36 7362 -2
rect 6970 -74 7362 -36
rect 6970 -108 6988 -74
rect 7022 -108 7310 -74
rect 7344 -108 7362 -74
rect 6970 -128 7362 -108
rect 7614 286 8006 306
rect 7614 252 7632 286
rect 7666 252 7954 286
rect 7988 252 8006 286
rect 7614 214 8006 252
rect 7614 180 7632 214
rect 7666 180 7954 214
rect 7988 180 8006 214
rect 7614 142 8006 180
rect 7614 108 7632 142
rect 7666 108 7954 142
rect 7988 108 8006 142
rect 7614 70 8006 108
rect 7614 36 7632 70
rect 7666 36 7954 70
rect 7988 36 8006 70
rect 7614 -2 8006 36
rect 7614 -36 7632 -2
rect 7666 -36 7954 -2
rect 7988 -36 8006 -2
rect 7614 -74 8006 -36
rect 7614 -108 7632 -74
rect 7666 -108 7954 -74
rect 7988 -108 8006 -74
rect 7614 -128 8006 -108
rect 0 -429 222 -395
rect 256 -429 276 -395
rect 0 -467 276 -429
rect 0 -501 222 -467
rect 256 -501 276 -467
rect 0 -539 276 -501
rect 0 -573 222 -539
rect 256 -573 276 -539
rect 0 -611 276 -573
rect 0 -645 222 -611
rect 256 -645 276 -611
rect 0 -683 276 -645
rect 0 -717 222 -683
rect 256 -717 276 -683
rect 0 -755 276 -717
rect 0 -789 222 -755
rect 256 -789 276 -755
rect 0 -812 276 -789
rect 526 -395 918 -374
rect 526 -429 544 -395
rect 578 -429 866 -395
rect 900 -429 918 -395
rect 526 -467 918 -429
rect 526 -501 544 -467
rect 578 -501 866 -467
rect 900 -501 918 -467
rect 526 -539 918 -501
rect 526 -573 544 -539
rect 578 -573 866 -539
rect 900 -573 918 -539
rect 526 -611 918 -573
rect 526 -645 544 -611
rect 578 -645 866 -611
rect 900 -645 918 -611
rect 526 -683 918 -645
rect 526 -717 544 -683
rect 578 -717 866 -683
rect 900 -717 918 -683
rect 526 -755 918 -717
rect 526 -789 544 -755
rect 578 -789 866 -755
rect 900 -789 918 -755
rect 526 -808 918 -789
rect 1170 -395 1562 -374
rect 1170 -429 1188 -395
rect 1222 -429 1510 -395
rect 1544 -429 1562 -395
rect 1170 -467 1562 -429
rect 1170 -501 1188 -467
rect 1222 -501 1510 -467
rect 1544 -501 1562 -467
rect 1170 -539 1562 -501
rect 1170 -573 1188 -539
rect 1222 -573 1510 -539
rect 1544 -573 1562 -539
rect 1170 -611 1562 -573
rect 1170 -645 1188 -611
rect 1222 -645 1510 -611
rect 1544 -645 1562 -611
rect 1170 -683 1562 -645
rect 1170 -717 1188 -683
rect 1222 -717 1510 -683
rect 1544 -717 1562 -683
rect 1170 -755 1562 -717
rect 1170 -789 1188 -755
rect 1222 -789 1510 -755
rect 1544 -789 1562 -755
rect 1170 -808 1562 -789
rect 1814 -395 2206 -374
rect 1814 -429 1832 -395
rect 1866 -429 2154 -395
rect 2188 -429 2206 -395
rect 1814 -467 2206 -429
rect 1814 -501 1832 -467
rect 1866 -501 2154 -467
rect 2188 -501 2206 -467
rect 1814 -539 2206 -501
rect 1814 -573 1832 -539
rect 1866 -573 2154 -539
rect 2188 -573 2206 -539
rect 1814 -611 2206 -573
rect 1814 -645 1832 -611
rect 1866 -645 2154 -611
rect 2188 -645 2206 -611
rect 1814 -683 2206 -645
rect 1814 -717 1832 -683
rect 1866 -717 2154 -683
rect 2188 -717 2206 -683
rect 1814 -755 2206 -717
rect 1814 -789 1832 -755
rect 1866 -789 2154 -755
rect 2188 -789 2206 -755
rect 1814 -808 2206 -789
rect 2458 -395 2850 -374
rect 2458 -429 2476 -395
rect 2510 -429 2798 -395
rect 2832 -429 2850 -395
rect 2458 -467 2850 -429
rect 2458 -501 2476 -467
rect 2510 -501 2798 -467
rect 2832 -501 2850 -467
rect 2458 -539 2850 -501
rect 2458 -573 2476 -539
rect 2510 -573 2798 -539
rect 2832 -573 2850 -539
rect 2458 -611 2850 -573
rect 2458 -645 2476 -611
rect 2510 -645 2798 -611
rect 2832 -645 2850 -611
rect 2458 -683 2850 -645
rect 2458 -717 2476 -683
rect 2510 -717 2798 -683
rect 2832 -717 2850 -683
rect 2458 -755 2850 -717
rect 2458 -789 2476 -755
rect 2510 -789 2798 -755
rect 2832 -789 2850 -755
rect 2458 -808 2850 -789
rect 3106 -395 3490 -382
rect 3106 -429 3120 -395
rect 3154 -429 3442 -395
rect 3476 -429 3490 -395
rect 3106 -467 3490 -429
rect 3106 -501 3120 -467
rect 3154 -501 3442 -467
rect 3476 -501 3490 -467
rect 3106 -539 3490 -501
rect 3106 -573 3120 -539
rect 3154 -573 3442 -539
rect 3476 -573 3490 -539
rect 3106 -611 3490 -573
rect 3106 -645 3120 -611
rect 3154 -645 3442 -611
rect 3476 -645 3490 -611
rect 3106 -683 3490 -645
rect 3106 -717 3120 -683
rect 3154 -717 3442 -683
rect 3476 -717 3490 -683
rect 3106 -755 3490 -717
rect 3106 -789 3120 -755
rect 3154 -789 3442 -755
rect 3476 -789 3490 -755
rect 3106 -804 3490 -789
rect 3750 -395 4134 -378
rect 3750 -429 3764 -395
rect 3798 -429 4086 -395
rect 4120 -429 4134 -395
rect 3750 -467 4134 -429
rect 3750 -501 3764 -467
rect 3798 -501 4086 -467
rect 4120 -501 4134 -467
rect 3750 -539 4134 -501
rect 3750 -573 3764 -539
rect 3798 -573 4086 -539
rect 4120 -573 4134 -539
rect 3750 -611 4134 -573
rect 3750 -645 3764 -611
rect 3798 -645 4086 -611
rect 4120 -645 4134 -611
rect 3750 -683 4134 -645
rect 3750 -717 3764 -683
rect 3798 -717 4086 -683
rect 4120 -717 4134 -683
rect 3750 -755 4134 -717
rect 3750 -789 3764 -755
rect 3798 -789 4086 -755
rect 4120 -789 4134 -755
rect 3750 -800 4134 -789
rect 4390 -395 4782 -374
rect 4390 -429 4408 -395
rect 4442 -429 4730 -395
rect 4764 -429 4782 -395
rect 4390 -467 4782 -429
rect 4390 -501 4408 -467
rect 4442 -501 4730 -467
rect 4764 -501 4782 -467
rect 4390 -539 4782 -501
rect 4390 -573 4408 -539
rect 4442 -573 4730 -539
rect 4764 -573 4782 -539
rect 4390 -611 4782 -573
rect 4390 -645 4408 -611
rect 4442 -645 4730 -611
rect 4764 -645 4782 -611
rect 4390 -683 4782 -645
rect 4390 -717 4408 -683
rect 4442 -717 4730 -683
rect 4764 -717 4782 -683
rect 4390 -755 4782 -717
rect 4390 -789 4408 -755
rect 4442 -789 4730 -755
rect 4764 -789 4782 -755
rect 4390 -808 4782 -789
rect 5034 -395 5426 -374
rect 5034 -429 5052 -395
rect 5086 -429 5374 -395
rect 5408 -429 5426 -395
rect 5034 -467 5426 -429
rect 5034 -501 5052 -467
rect 5086 -501 5374 -467
rect 5408 -501 5426 -467
rect 5034 -539 5426 -501
rect 5034 -573 5052 -539
rect 5086 -573 5374 -539
rect 5408 -573 5426 -539
rect 5034 -611 5426 -573
rect 5034 -645 5052 -611
rect 5086 -645 5374 -611
rect 5408 -645 5426 -611
rect 5034 -683 5426 -645
rect 5034 -717 5052 -683
rect 5086 -717 5374 -683
rect 5408 -717 5426 -683
rect 5034 -755 5426 -717
rect 5034 -789 5052 -755
rect 5086 -789 5374 -755
rect 5408 -789 5426 -755
rect 5034 -808 5426 -789
rect 5678 -395 6070 -374
rect 5678 -429 5696 -395
rect 5730 -429 6018 -395
rect 6052 -429 6070 -395
rect 5678 -467 6070 -429
rect 5678 -501 5696 -467
rect 5730 -501 6018 -467
rect 6052 -501 6070 -467
rect 5678 -539 6070 -501
rect 5678 -573 5696 -539
rect 5730 -573 6018 -539
rect 6052 -573 6070 -539
rect 5678 -611 6070 -573
rect 5678 -645 5696 -611
rect 5730 -645 6018 -611
rect 6052 -645 6070 -611
rect 5678 -683 6070 -645
rect 5678 -717 5696 -683
rect 5730 -717 6018 -683
rect 6052 -717 6070 -683
rect 5678 -755 6070 -717
rect 5678 -789 5696 -755
rect 5730 -789 6018 -755
rect 6052 -789 6070 -755
rect 5678 -808 6070 -789
rect 6322 -395 6714 -374
rect 6322 -429 6340 -395
rect 6374 -429 6662 -395
rect 6696 -429 6714 -395
rect 6322 -467 6714 -429
rect 6322 -501 6340 -467
rect 6374 -501 6662 -467
rect 6696 -501 6714 -467
rect 6322 -539 6714 -501
rect 6322 -573 6340 -539
rect 6374 -573 6662 -539
rect 6696 -573 6714 -539
rect 6322 -611 6714 -573
rect 6322 -645 6340 -611
rect 6374 -645 6662 -611
rect 6696 -645 6714 -611
rect 6322 -683 6714 -645
rect 6322 -717 6340 -683
rect 6374 -717 6662 -683
rect 6696 -717 6714 -683
rect 6322 -755 6714 -717
rect 6322 -789 6340 -755
rect 6374 -789 6662 -755
rect 6696 -789 6714 -755
rect 6322 -808 6714 -789
rect 6968 -395 7354 -380
rect 6968 -429 6984 -395
rect 7018 -429 7306 -395
rect 7340 -429 7354 -395
rect 6968 -467 7354 -429
rect 6968 -501 6984 -467
rect 7018 -501 7306 -467
rect 7340 -501 7354 -467
rect 6968 -539 7354 -501
rect 6968 -573 6984 -539
rect 7018 -573 7306 -539
rect 7340 -573 7354 -539
rect 6968 -611 7354 -573
rect 6968 -645 6984 -611
rect 7018 -645 7306 -611
rect 7340 -645 7354 -611
rect 6968 -683 7354 -645
rect 6968 -717 6984 -683
rect 7018 -717 7306 -683
rect 7340 -717 7354 -683
rect 6968 -755 7354 -717
rect 6968 -789 6984 -755
rect 7018 -789 7306 -755
rect 7340 -789 7354 -755
rect 6968 -804 7354 -789
rect 7610 -395 8002 -374
rect 7610 -429 7628 -395
rect 7662 -429 7950 -395
rect 7984 -429 8002 -395
rect 7610 -467 8002 -429
rect 7610 -501 7628 -467
rect 7662 -501 7950 -467
rect 7984 -501 8002 -467
rect 7610 -539 8002 -501
rect 7610 -573 7628 -539
rect 7662 -573 7950 -539
rect 7984 -573 8002 -539
rect 7610 -611 8002 -573
rect 7610 -645 7628 -611
rect 7662 -645 7950 -611
rect 7984 -645 8002 -611
rect 7610 -683 8002 -645
rect 7610 -717 7628 -683
rect 7662 -717 7950 -683
rect 7984 -717 8002 -683
rect 7610 -755 8002 -717
rect 7610 -789 7628 -755
rect 7662 -789 7950 -755
rect 7984 -789 8002 -755
rect 7610 -808 8002 -789
rect 204 -2202 596 -2182
rect 204 -2236 222 -2202
rect 256 -2236 544 -2202
rect 578 -2236 596 -2202
rect 204 -2274 596 -2236
rect 204 -2308 222 -2274
rect 256 -2308 544 -2274
rect 578 -2308 596 -2274
rect 204 -2346 596 -2308
rect 204 -2380 222 -2346
rect 256 -2380 544 -2346
rect 578 -2380 596 -2346
rect 204 -2418 596 -2380
rect 204 -2452 222 -2418
rect 256 -2452 544 -2418
rect 578 -2452 596 -2418
rect 204 -2490 596 -2452
rect 204 -2524 222 -2490
rect 256 -2524 544 -2490
rect 578 -2524 596 -2490
rect 204 -2562 596 -2524
rect 204 -2596 222 -2562
rect 256 -2596 544 -2562
rect 578 -2596 596 -2562
rect 204 -2616 596 -2596
rect 848 -2202 1240 -2182
rect 848 -2236 866 -2202
rect 900 -2236 1188 -2202
rect 1222 -2236 1240 -2202
rect 848 -2274 1240 -2236
rect 848 -2308 866 -2274
rect 900 -2308 1188 -2274
rect 1222 -2308 1240 -2274
rect 848 -2346 1240 -2308
rect 848 -2380 866 -2346
rect 900 -2380 1188 -2346
rect 1222 -2380 1240 -2346
rect 848 -2418 1240 -2380
rect 848 -2452 866 -2418
rect 900 -2452 1188 -2418
rect 1222 -2452 1240 -2418
rect 848 -2490 1240 -2452
rect 848 -2524 866 -2490
rect 900 -2524 1188 -2490
rect 1222 -2524 1240 -2490
rect 848 -2562 1240 -2524
rect 848 -2596 866 -2562
rect 900 -2596 1188 -2562
rect 1222 -2596 1240 -2562
rect 848 -2616 1240 -2596
rect 1492 -2202 1884 -2182
rect 1492 -2236 1510 -2202
rect 1544 -2236 1832 -2202
rect 1866 -2236 1884 -2202
rect 1492 -2274 1884 -2236
rect 1492 -2308 1510 -2274
rect 1544 -2308 1832 -2274
rect 1866 -2308 1884 -2274
rect 1492 -2346 1884 -2308
rect 1492 -2380 1510 -2346
rect 1544 -2380 1832 -2346
rect 1866 -2380 1884 -2346
rect 1492 -2418 1884 -2380
rect 1492 -2452 1510 -2418
rect 1544 -2452 1832 -2418
rect 1866 -2452 1884 -2418
rect 1492 -2490 1884 -2452
rect 1492 -2524 1510 -2490
rect 1544 -2524 1832 -2490
rect 1866 -2524 1884 -2490
rect 1492 -2562 1884 -2524
rect 1492 -2596 1510 -2562
rect 1544 -2596 1832 -2562
rect 1866 -2596 1884 -2562
rect 1492 -2616 1884 -2596
rect 2136 -2202 2528 -2182
rect 2136 -2236 2154 -2202
rect 2188 -2236 2476 -2202
rect 2510 -2236 2528 -2202
rect 2136 -2274 2528 -2236
rect 2136 -2308 2154 -2274
rect 2188 -2308 2476 -2274
rect 2510 -2308 2528 -2274
rect 2136 -2346 2528 -2308
rect 2136 -2380 2154 -2346
rect 2188 -2380 2476 -2346
rect 2510 -2380 2528 -2346
rect 2136 -2418 2528 -2380
rect 2136 -2452 2154 -2418
rect 2188 -2452 2476 -2418
rect 2510 -2452 2528 -2418
rect 2136 -2490 2528 -2452
rect 2136 -2524 2154 -2490
rect 2188 -2524 2476 -2490
rect 2510 -2524 2528 -2490
rect 2136 -2562 2528 -2524
rect 2136 -2596 2154 -2562
rect 2188 -2596 2476 -2562
rect 2510 -2596 2528 -2562
rect 2136 -2616 2528 -2596
rect 2780 -2202 3172 -2182
rect 2780 -2236 2798 -2202
rect 2832 -2236 3120 -2202
rect 3154 -2236 3172 -2202
rect 2780 -2274 3172 -2236
rect 2780 -2308 2798 -2274
rect 2832 -2308 3120 -2274
rect 3154 -2308 3172 -2274
rect 2780 -2346 3172 -2308
rect 2780 -2380 2798 -2346
rect 2832 -2380 3120 -2346
rect 3154 -2380 3172 -2346
rect 2780 -2418 3172 -2380
rect 2780 -2452 2798 -2418
rect 2832 -2452 3120 -2418
rect 3154 -2452 3172 -2418
rect 2780 -2490 3172 -2452
rect 2780 -2524 2798 -2490
rect 2832 -2524 3120 -2490
rect 3154 -2524 3172 -2490
rect 2780 -2562 3172 -2524
rect 2780 -2596 2798 -2562
rect 2832 -2596 3120 -2562
rect 3154 -2596 3172 -2562
rect 2780 -2616 3172 -2596
rect 3424 -2202 3816 -2182
rect 3424 -2236 3442 -2202
rect 3476 -2236 3764 -2202
rect 3798 -2236 3816 -2202
rect 3424 -2274 3816 -2236
rect 3424 -2308 3442 -2274
rect 3476 -2308 3764 -2274
rect 3798 -2308 3816 -2274
rect 3424 -2346 3816 -2308
rect 3424 -2380 3442 -2346
rect 3476 -2380 3764 -2346
rect 3798 -2380 3816 -2346
rect 3424 -2418 3816 -2380
rect 3424 -2452 3442 -2418
rect 3476 -2452 3764 -2418
rect 3798 -2452 3816 -2418
rect 3424 -2490 3816 -2452
rect 3424 -2524 3442 -2490
rect 3476 -2524 3764 -2490
rect 3798 -2524 3816 -2490
rect 3424 -2562 3816 -2524
rect 3424 -2596 3442 -2562
rect 3476 -2596 3764 -2562
rect 3798 -2596 3816 -2562
rect 3424 -2616 3816 -2596
rect 4068 -2202 4460 -2182
rect 4068 -2236 4086 -2202
rect 4120 -2236 4408 -2202
rect 4442 -2236 4460 -2202
rect 4068 -2274 4460 -2236
rect 4068 -2308 4086 -2274
rect 4120 -2308 4408 -2274
rect 4442 -2308 4460 -2274
rect 4068 -2346 4460 -2308
rect 4068 -2380 4086 -2346
rect 4120 -2380 4408 -2346
rect 4442 -2380 4460 -2346
rect 4068 -2418 4460 -2380
rect 4068 -2452 4086 -2418
rect 4120 -2452 4408 -2418
rect 4442 -2452 4460 -2418
rect 4068 -2490 4460 -2452
rect 4068 -2524 4086 -2490
rect 4120 -2524 4408 -2490
rect 4442 -2524 4460 -2490
rect 4068 -2562 4460 -2524
rect 4068 -2596 4086 -2562
rect 4120 -2596 4408 -2562
rect 4442 -2596 4460 -2562
rect 4068 -2616 4460 -2596
rect 4712 -2202 5104 -2182
rect 4712 -2236 4730 -2202
rect 4764 -2236 5052 -2202
rect 5086 -2236 5104 -2202
rect 4712 -2274 5104 -2236
rect 4712 -2308 4730 -2274
rect 4764 -2308 5052 -2274
rect 5086 -2308 5104 -2274
rect 4712 -2346 5104 -2308
rect 4712 -2380 4730 -2346
rect 4764 -2380 5052 -2346
rect 5086 -2380 5104 -2346
rect 4712 -2418 5104 -2380
rect 4712 -2452 4730 -2418
rect 4764 -2452 5052 -2418
rect 5086 -2452 5104 -2418
rect 4712 -2490 5104 -2452
rect 4712 -2524 4730 -2490
rect 4764 -2524 5052 -2490
rect 5086 -2524 5104 -2490
rect 4712 -2562 5104 -2524
rect 4712 -2596 4730 -2562
rect 4764 -2596 5052 -2562
rect 5086 -2596 5104 -2562
rect 4712 -2616 5104 -2596
rect 5356 -2202 5748 -2182
rect 5356 -2236 5374 -2202
rect 5408 -2236 5696 -2202
rect 5730 -2236 5748 -2202
rect 5356 -2274 5748 -2236
rect 5356 -2308 5374 -2274
rect 5408 -2308 5696 -2274
rect 5730 -2308 5748 -2274
rect 5356 -2346 5748 -2308
rect 5356 -2380 5374 -2346
rect 5408 -2380 5696 -2346
rect 5730 -2380 5748 -2346
rect 5356 -2418 5748 -2380
rect 5356 -2452 5374 -2418
rect 5408 -2452 5696 -2418
rect 5730 -2452 5748 -2418
rect 5356 -2490 5748 -2452
rect 5356 -2524 5374 -2490
rect 5408 -2524 5696 -2490
rect 5730 -2524 5748 -2490
rect 5356 -2562 5748 -2524
rect 5356 -2596 5374 -2562
rect 5408 -2596 5696 -2562
rect 5730 -2596 5748 -2562
rect 5356 -2616 5748 -2596
rect 6000 -2202 6392 -2182
rect 6000 -2236 6018 -2202
rect 6052 -2236 6340 -2202
rect 6374 -2236 6392 -2202
rect 6000 -2274 6392 -2236
rect 6000 -2308 6018 -2274
rect 6052 -2308 6340 -2274
rect 6374 -2308 6392 -2274
rect 6000 -2346 6392 -2308
rect 6000 -2380 6018 -2346
rect 6052 -2380 6340 -2346
rect 6374 -2380 6392 -2346
rect 6000 -2418 6392 -2380
rect 6000 -2452 6018 -2418
rect 6052 -2452 6340 -2418
rect 6374 -2452 6392 -2418
rect 6000 -2490 6392 -2452
rect 6000 -2524 6018 -2490
rect 6052 -2524 6340 -2490
rect 6374 -2524 6392 -2490
rect 6000 -2562 6392 -2524
rect 6000 -2596 6018 -2562
rect 6052 -2596 6340 -2562
rect 6374 -2596 6392 -2562
rect 6000 -2616 6392 -2596
rect 6644 -2202 7036 -2182
rect 6644 -2236 6662 -2202
rect 6696 -2236 6984 -2202
rect 7018 -2236 7036 -2202
rect 6644 -2274 7036 -2236
rect 6644 -2308 6662 -2274
rect 6696 -2308 6984 -2274
rect 7018 -2308 7036 -2274
rect 6644 -2346 7036 -2308
rect 6644 -2380 6662 -2346
rect 6696 -2380 6984 -2346
rect 7018 -2380 7036 -2346
rect 6644 -2418 7036 -2380
rect 6644 -2452 6662 -2418
rect 6696 -2452 6984 -2418
rect 7018 -2452 7036 -2418
rect 6644 -2490 7036 -2452
rect 6644 -2524 6662 -2490
rect 6696 -2524 6984 -2490
rect 7018 -2524 7036 -2490
rect 6644 -2562 7036 -2524
rect 6644 -2596 6662 -2562
rect 6696 -2596 6984 -2562
rect 7018 -2596 7036 -2562
rect 6644 -2616 7036 -2596
rect 7288 -2202 7680 -2182
rect 7288 -2236 7306 -2202
rect 7340 -2236 7628 -2202
rect 7662 -2236 7680 -2202
rect 7288 -2274 7680 -2236
rect 7288 -2308 7306 -2274
rect 7340 -2308 7628 -2274
rect 7662 -2308 7680 -2274
rect 7288 -2346 7680 -2308
rect 7288 -2380 7306 -2346
rect 7340 -2380 7628 -2346
rect 7662 -2380 7680 -2346
rect 7288 -2418 7680 -2380
rect 7288 -2452 7306 -2418
rect 7340 -2452 7628 -2418
rect 7662 -2452 7680 -2418
rect 7288 -2490 7680 -2452
rect 7288 -2524 7306 -2490
rect 7340 -2524 7628 -2490
rect 7662 -2524 7680 -2490
rect 7288 -2562 7680 -2524
rect 7288 -2596 7306 -2562
rect 7340 -2596 7628 -2562
rect 7662 -2596 7680 -2562
rect 7288 -2616 7680 -2596
rect 7936 -2202 8002 -2182
rect 7936 -2236 7950 -2202
rect 7984 -2236 8002 -2202
rect 7936 -2274 8002 -2236
rect 7936 -2308 7950 -2274
rect 7984 -2308 8002 -2274
rect 7936 -2346 8002 -2308
rect 7936 -2380 7950 -2346
rect 7984 -2380 8002 -2346
rect 7936 -2418 8002 -2380
rect 7936 -2452 7950 -2418
rect 7984 -2452 8002 -2418
rect 7936 -2490 8002 -2452
rect 7936 -2524 7950 -2490
rect 7984 -2524 8002 -2490
rect 7936 -2562 8002 -2524
rect 7936 -2596 7950 -2562
rect 7984 -2596 8002 -2562
rect 7936 -2756 8002 -2596
rect 7192 -2813 8012 -2756
rect 7192 -2929 7256 -2813
rect 7948 -2929 8012 -2813
rect 7192 -2982 8012 -2929
<< via1 >>
rect 7267 2329 7959 2509
rect 7256 -2929 7948 -2813
<< metal2 >>
rect 7222 2509 8004 2532
rect 7222 2329 7267 2509
rect 7959 2329 8004 2509
rect 7222 2308 8004 2329
rect 7196 -2813 8006 -2760
rect 7196 -2929 7256 -2813
rect 7948 -2929 8006 -2813
rect 7196 -2992 8006 -2929
<< labels >>
rlabel metal1 s 8 -804 196 296 4 vcm
port 1 nsew
rlabel metal2 s 7212 -2982 7996 -2772 4 GND
port 2 nsew
rlabel locali s 432 -272 7976 -228 4 GND
port 2 nsew
rlabel metal2 s 7236 2316 7992 2520 4 VDD
port 3 nsew
<< end >>
