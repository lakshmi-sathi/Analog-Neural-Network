magic
tech sky130A
magscale 1 2
timestamp 1627668659
<< error_p >>
rect -29 592 29 598
rect -29 558 -17 592
rect -29 552 29 558
rect -29 -558 29 -552
rect -29 -592 -17 -558
rect -29 -598 29 -592
<< pwell >>
rect -211 -730 211 730
<< nmos >>
rect -15 -520 15 520
<< ndiff >>
rect -73 508 -15 520
rect -73 -508 -61 508
rect -27 -508 -15 508
rect -73 -520 -15 -508
rect 15 508 73 520
rect 15 -508 27 508
rect 61 -508 73 508
rect 15 -520 73 -508
<< ndiffc >>
rect -61 -508 -27 508
rect 27 -508 61 508
<< psubdiff >>
rect -175 660 -79 694
rect 79 660 175 694
rect -175 598 -141 660
rect 141 598 175 660
rect -175 -660 -141 -598
rect 141 -660 175 -598
rect -175 -694 -79 -660
rect 79 -694 175 -660
<< psubdiffcont >>
rect -79 660 79 694
rect -175 -598 -141 598
rect 141 -598 175 598
rect -79 -694 79 -660
<< poly >>
rect -33 592 33 608
rect -33 558 -17 592
rect 17 558 33 592
rect -33 542 33 558
rect -15 520 15 542
rect -15 -542 15 -520
rect -33 -558 33 -542
rect -33 -592 -17 -558
rect 17 -592 33 -558
rect -33 -608 33 -592
<< polycont >>
rect -17 558 17 592
rect -17 -592 17 -558
<< locali >>
rect -175 660 -79 694
rect 79 660 175 694
rect -175 598 -141 660
rect 141 598 175 660
rect -33 558 -17 592
rect 17 558 33 592
rect -61 508 -27 524
rect -61 -524 -27 -508
rect 27 508 61 524
rect 27 -524 61 -508
rect -33 -592 -17 -558
rect 17 -592 33 -558
rect -175 -660 -141 -598
rect 141 -660 175 -598
rect -175 -694 -79 -660
rect 79 -694 175 -660
<< viali >>
rect -17 558 17 592
rect -61 -508 -27 508
rect 27 -508 61 508
rect -17 -592 17 -558
<< metal1 >>
rect -29 592 29 598
rect -29 558 -17 592
rect 17 558 29 592
rect -29 552 29 558
rect -67 508 -21 520
rect -67 -508 -61 508
rect -27 -508 -21 508
rect -67 -520 -21 -508
rect 21 508 67 520
rect 21 -508 27 508
rect 61 -508 67 508
rect 21 -520 67 -508
rect -29 -558 29 -552
rect -29 -592 -17 -558
rect 17 -592 29 -558
rect -29 -598 29 -592
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -677 158 677
string parameters w 5.2 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
