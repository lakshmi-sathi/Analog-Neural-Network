magic
tech sky130A
magscale 1 2
timestamp 1627926120
<< xpolycontact >>
rect -35 638 35 1070
rect -35 -1070 35 -638
<< xpolyres >>
rect -35 -638 35 638
<< viali >>
rect -17 1016 17 1050
rect -17 944 17 978
rect -17 872 17 906
rect -17 800 17 834
rect -17 728 17 762
rect -17 656 17 690
rect -17 -691 17 -657
rect -17 -763 17 -729
rect -17 -835 17 -801
rect -17 -907 17 -873
rect -17 -979 17 -945
rect -17 -1051 17 -1017
<< metal1 >>
rect -25 1050 25 1064
rect -25 1016 -17 1050
rect 17 1016 25 1050
rect -25 978 25 1016
rect -25 944 -17 978
rect 17 944 25 978
rect -25 906 25 944
rect -25 872 -17 906
rect 17 872 25 906
rect -25 834 25 872
rect -25 800 -17 834
rect 17 800 25 834
rect -25 762 25 800
rect -25 728 -17 762
rect 17 728 25 762
rect -25 690 25 728
rect -25 656 -17 690
rect 17 656 25 690
rect -25 643 25 656
rect -25 -657 25 -643
rect -25 -691 -17 -657
rect 17 -691 25 -657
rect -25 -729 25 -691
rect -25 -763 -17 -729
rect 17 -763 25 -729
rect -25 -801 25 -763
rect -25 -835 -17 -801
rect 17 -835 25 -801
rect -25 -873 25 -835
rect -25 -907 -17 -873
rect 17 -907 25 -873
rect -25 -945 25 -907
rect -25 -979 -17 -945
rect 17 -979 25 -945
rect -25 -1017 25 -979
rect -25 -1051 -17 -1017
rect 17 -1051 25 -1017
rect -25 -1064 25 -1051
<< end >>
