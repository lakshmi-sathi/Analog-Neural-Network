magic
tech sky130A
magscale 1 2
timestamp 1627883883
<< psubdiff >>
rect 408 -272 432 -228
rect 7976 -272 8000 -228
<< psubdiffcont >>
rect 432 -272 7976 -228
<< xpolycontact >>
rect 208 1681 278 2113
rect 208 -127 278 305
rect 530 1681 600 2113
rect 530 -127 600 305
rect 852 1681 922 2113
rect 852 -127 922 305
rect 1174 1681 1244 2113
rect 1174 -127 1244 305
rect 1496 1681 1566 2113
rect 1496 -127 1566 305
rect 1818 1681 1888 2113
rect 1818 -127 1888 305
rect 2140 1681 2210 2113
rect 2140 -127 2210 305
rect 2462 1681 2532 2113
rect 2462 -127 2532 305
rect 2784 1681 2854 2113
rect 2784 -127 2854 305
rect 3106 1681 3176 2113
rect 3106 -127 3176 305
rect 3428 1681 3498 2113
rect 3428 -127 3498 305
rect 3750 1681 3820 2113
rect 3750 -127 3820 305
rect 4072 1681 4142 2113
rect 4072 -127 4142 305
rect 4394 1681 4464 2113
rect 4394 -127 4464 305
rect 4716 1681 4786 2113
rect 4716 -127 4786 305
rect 5038 1681 5108 2113
rect 5038 -127 5108 305
rect 5360 1681 5430 2113
rect 5360 -127 5430 305
rect 5682 1681 5752 2113
rect 5682 -127 5752 305
rect 6004 1681 6074 2113
rect 6004 -127 6074 305
rect 6326 1681 6396 2113
rect 6326 -127 6396 305
rect 6648 1681 6718 2113
rect 6648 -127 6718 305
rect 6970 1681 7040 2113
rect 6970 -127 7040 305
rect 7292 1681 7362 2113
rect 7292 -127 7362 305
rect 7614 1681 7684 2113
rect 7614 -127 7684 305
rect 7936 1681 8006 2113
rect 7936 -127 8006 305
rect 204 -807 274 -375
rect 204 -2615 274 -2183
rect 526 -807 596 -375
rect 526 -2615 596 -2183
rect 848 -807 918 -375
rect 848 -2615 918 -2183
rect 1170 -807 1240 -375
rect 1170 -2615 1240 -2183
rect 1492 -807 1562 -375
rect 1492 -2615 1562 -2183
rect 1814 -807 1884 -375
rect 1814 -2615 1884 -2183
rect 2136 -807 2206 -375
rect 2136 -2615 2206 -2183
rect 2458 -807 2528 -375
rect 2458 -2615 2528 -2183
rect 2780 -807 2850 -375
rect 2780 -2615 2850 -2183
rect 3102 -807 3172 -375
rect 3102 -2615 3172 -2183
rect 3424 -807 3494 -375
rect 3424 -2615 3494 -2183
rect 3746 -807 3816 -375
rect 3746 -2615 3816 -2183
rect 4068 -807 4138 -375
rect 4068 -2615 4138 -2183
rect 4390 -807 4460 -375
rect 4390 -2615 4460 -2183
rect 4712 -807 4782 -375
rect 4712 -2615 4782 -2183
rect 5034 -807 5104 -375
rect 5034 -2615 5104 -2183
rect 5356 -807 5426 -375
rect 5356 -2615 5426 -2183
rect 5678 -807 5748 -375
rect 5678 -2615 5748 -2183
rect 6000 -807 6070 -375
rect 6000 -2615 6070 -2183
rect 6322 -807 6392 -375
rect 6322 -2615 6392 -2183
rect 6644 -807 6714 -375
rect 6644 -2615 6714 -2183
rect 6966 -807 7036 -375
rect 6966 -2615 7036 -2183
rect 7288 -807 7358 -375
rect 7288 -2615 7358 -2183
rect 7610 -807 7680 -375
rect 7610 -2615 7680 -2183
rect 7932 -807 8002 -375
rect 7932 -2615 8002 -2183
<< xpolyres >>
rect 208 305 278 1681
rect 530 305 600 1681
rect 852 305 922 1681
rect 1174 305 1244 1681
rect 1496 305 1566 1681
rect 1818 305 1888 1681
rect 2140 305 2210 1681
rect 2462 305 2532 1681
rect 2784 305 2854 1681
rect 3106 305 3176 1681
rect 3428 305 3498 1681
rect 3750 305 3820 1681
rect 4072 305 4142 1681
rect 4394 305 4464 1681
rect 4716 305 4786 1681
rect 5038 305 5108 1681
rect 5360 305 5430 1681
rect 5682 305 5752 1681
rect 6004 305 6074 1681
rect 6326 305 6396 1681
rect 6648 305 6718 1681
rect 6970 305 7040 1681
rect 7292 305 7362 1681
rect 7614 305 7684 1681
rect 7936 305 8006 1681
rect 204 -2183 274 -807
rect 526 -2183 596 -807
rect 848 -2183 918 -807
rect 1170 -2183 1240 -807
rect 1492 -2183 1562 -807
rect 1814 -2183 1884 -807
rect 2136 -2183 2206 -807
rect 2458 -2183 2528 -807
rect 2780 -2183 2850 -807
rect 3102 -2183 3172 -807
rect 3424 -2183 3494 -807
rect 3746 -2183 3816 -807
rect 4068 -2183 4138 -807
rect 4390 -2183 4460 -807
rect 4712 -2183 4782 -807
rect 5034 -2183 5104 -807
rect 5356 -2183 5426 -807
rect 5678 -2183 5748 -807
rect 6000 -2183 6070 -807
rect 6322 -2183 6392 -807
rect 6644 -2183 6714 -807
rect 6966 -2183 7036 -807
rect 7288 -2183 7358 -807
rect 7610 -2183 7680 -807
rect 7932 -2183 8002 -807
<< locali >>
rect 416 -272 432 -228
rect 7976 -272 7992 -228
<< viali >>
rect 224 1698 262 2095
rect 546 1698 584 2095
rect 868 1698 906 2095
rect 1190 1698 1228 2095
rect 1512 1698 1550 2095
rect 1834 1698 1872 2095
rect 2156 1698 2194 2095
rect 2478 1698 2516 2095
rect 2800 1698 2838 2095
rect 3122 1698 3160 2095
rect 3444 1698 3482 2095
rect 3766 1698 3804 2095
rect 4088 1698 4126 2095
rect 4410 1698 4448 2095
rect 4732 1698 4770 2095
rect 5054 1698 5092 2095
rect 5376 1698 5414 2095
rect 5698 1698 5736 2095
rect 6020 1698 6058 2095
rect 6342 1698 6380 2095
rect 6664 1698 6702 2095
rect 6986 1698 7024 2095
rect 7308 1698 7346 2095
rect 7630 1698 7668 2095
rect 7952 1698 7990 2095
rect 224 -109 262 288
rect 546 -109 584 288
rect 868 -109 906 288
rect 1190 -109 1228 288
rect 1512 -109 1550 288
rect 1834 -109 1872 288
rect 2156 -109 2194 288
rect 2478 -109 2516 288
rect 2800 -109 2838 288
rect 3122 -109 3160 288
rect 3444 -109 3482 288
rect 3766 -109 3804 288
rect 4088 -109 4126 288
rect 4410 -109 4448 288
rect 4732 -109 4770 288
rect 5054 -109 5092 288
rect 5376 -109 5414 288
rect 5698 -109 5736 288
rect 6020 -109 6058 288
rect 6342 -109 6380 288
rect 6664 -109 6702 288
rect 6986 -109 7024 288
rect 7308 -109 7346 288
rect 7630 -109 7668 288
rect 7952 -109 7990 288
rect 220 -790 258 -393
rect 542 -790 580 -393
rect 864 -790 902 -393
rect 1186 -790 1224 -393
rect 1508 -790 1546 -393
rect 1830 -790 1868 -393
rect 2152 -790 2190 -393
rect 2474 -790 2512 -393
rect 2796 -790 2834 -393
rect 3118 -790 3156 -393
rect 3440 -790 3478 -393
rect 3762 -790 3800 -393
rect 4084 -790 4122 -393
rect 4406 -790 4444 -393
rect 4728 -790 4766 -393
rect 5050 -790 5088 -393
rect 5372 -790 5410 -393
rect 5694 -790 5732 -393
rect 6016 -790 6054 -393
rect 6338 -790 6376 -393
rect 6660 -790 6698 -393
rect 6982 -790 7020 -393
rect 7304 -790 7342 -393
rect 7626 -790 7664 -393
rect 7948 -790 7986 -393
rect 220 -2597 258 -2200
rect 542 -2597 580 -2200
rect 864 -2597 902 -2200
rect 1186 -2597 1224 -2200
rect 1508 -2597 1546 -2200
rect 1830 -2597 1868 -2200
rect 2152 -2597 2190 -2200
rect 2474 -2597 2512 -2200
rect 2796 -2597 2834 -2200
rect 3118 -2597 3156 -2200
rect 3440 -2597 3478 -2200
rect 3762 -2597 3800 -2200
rect 4084 -2597 4122 -2200
rect 4406 -2597 4444 -2200
rect 4728 -2597 4766 -2200
rect 5050 -2597 5088 -2200
rect 5372 -2597 5410 -2200
rect 5694 -2597 5732 -2200
rect 6016 -2597 6054 -2200
rect 6338 -2597 6376 -2200
rect 6660 -2597 6698 -2200
rect 6982 -2597 7020 -2200
rect 7304 -2597 7342 -2200
rect 7626 -2597 7664 -2200
rect 7948 -2597 7986 -2200
<< metal1 >>
rect 7212 2512 8012 2542
rect 7212 2326 7252 2512
rect 7974 2326 8012 2512
rect 7212 2302 8012 2326
rect 208 2095 600 2114
rect 208 1698 224 2095
rect 262 1698 546 2095
rect 584 1698 600 2095
rect 208 1680 600 1698
rect 852 2095 1244 2114
rect 852 1698 868 2095
rect 906 1698 1190 2095
rect 1228 1698 1244 2095
rect 852 1680 1244 1698
rect 1496 2095 1888 2114
rect 1496 1698 1512 2095
rect 1550 1698 1834 2095
rect 1872 1698 1888 2095
rect 1496 1680 1888 1698
rect 2140 2095 2532 2114
rect 2140 1698 2156 2095
rect 2194 1698 2478 2095
rect 2516 1698 2532 2095
rect 2140 1680 2532 1698
rect 2784 2095 3176 2114
rect 2784 1698 2800 2095
rect 2838 1698 3122 2095
rect 3160 1698 3176 2095
rect 2784 1680 3176 1698
rect 3428 2095 3820 2114
rect 3428 1698 3444 2095
rect 3482 1698 3766 2095
rect 3804 1698 3820 2095
rect 3428 1680 3820 1698
rect 4072 2095 4464 2114
rect 4072 1698 4088 2095
rect 4126 1698 4410 2095
rect 4448 1698 4464 2095
rect 4072 1680 4464 1698
rect 4716 2095 5108 2114
rect 4716 1698 4732 2095
rect 4770 1698 5054 2095
rect 5092 1698 5108 2095
rect 4716 1680 5108 1698
rect 5360 2095 5752 2114
rect 5360 1698 5376 2095
rect 5414 1698 5698 2095
rect 5736 1698 5752 2095
rect 5360 1680 5752 1698
rect 6004 2095 6396 2114
rect 6004 1698 6020 2095
rect 6058 1698 6342 2095
rect 6380 1698 6396 2095
rect 6004 1680 6396 1698
rect 6648 2095 7040 2114
rect 6648 1698 6664 2095
rect 6702 1698 6986 2095
rect 7024 1698 7040 2095
rect 6648 1680 7040 1698
rect 7292 2095 7684 2114
rect 7292 1698 7308 2095
rect 7346 1698 7630 2095
rect 7668 1698 7684 2095
rect 7936 2095 8006 2302
rect 7936 2084 7952 2095
rect 7292 1680 7684 1698
rect 7946 1698 7952 2084
rect 7990 2084 8006 2095
rect 7990 1698 7996 2084
rect 7946 1686 7996 1698
rect 0 288 276 306
rect 0 -109 224 288
rect 262 -109 276 288
rect 0 -393 276 -109
rect 530 288 922 306
rect 530 -109 546 288
rect 584 -109 868 288
rect 906 -109 922 288
rect 530 -128 922 -109
rect 1174 288 1566 306
rect 1174 -109 1190 288
rect 1228 -109 1512 288
rect 1550 -109 1566 288
rect 1174 -128 1566 -109
rect 1818 288 2210 306
rect 1818 -109 1834 288
rect 1872 -109 2156 288
rect 2194 -109 2210 288
rect 1818 -128 2210 -109
rect 2462 288 2854 306
rect 2462 -109 2478 288
rect 2516 -109 2800 288
rect 2838 -109 2854 288
rect 2462 -128 2854 -109
rect 3106 288 3498 306
rect 3106 -109 3122 288
rect 3160 -109 3444 288
rect 3482 -109 3498 288
rect 3106 -128 3498 -109
rect 3750 288 4142 306
rect 3750 -109 3766 288
rect 3804 -109 4088 288
rect 4126 -109 4142 288
rect 3750 -128 4142 -109
rect 4394 288 4786 306
rect 4394 -109 4410 288
rect 4448 -109 4732 288
rect 4770 -109 4786 288
rect 4394 -128 4786 -109
rect 5038 288 5430 306
rect 5038 -109 5054 288
rect 5092 -109 5376 288
rect 5414 -109 5430 288
rect 5038 -128 5430 -109
rect 5682 288 6074 306
rect 5682 -109 5698 288
rect 5736 -109 6020 288
rect 6058 -109 6074 288
rect 5682 -128 6074 -109
rect 6326 288 6718 306
rect 6326 -109 6342 288
rect 6380 -109 6664 288
rect 6702 -109 6718 288
rect 6326 -128 6718 -109
rect 6970 288 7362 306
rect 6970 -109 6986 288
rect 7024 -109 7308 288
rect 7346 -109 7362 288
rect 6970 -128 7362 -109
rect 7614 288 8006 306
rect 7614 -109 7630 288
rect 7668 -109 7952 288
rect 7990 -109 8006 288
rect 7614 -128 8006 -109
rect 0 -790 220 -393
rect 258 -790 276 -393
rect 0 -812 276 -790
rect 526 -393 918 -374
rect 526 -790 542 -393
rect 580 -790 864 -393
rect 902 -790 918 -393
rect 526 -808 918 -790
rect 1170 -393 1562 -374
rect 1170 -790 1186 -393
rect 1224 -790 1508 -393
rect 1546 -790 1562 -393
rect 1170 -808 1562 -790
rect 1814 -393 2206 -374
rect 1814 -790 1830 -393
rect 1868 -790 2152 -393
rect 2190 -790 2206 -393
rect 1814 -808 2206 -790
rect 2458 -393 2850 -374
rect 2458 -790 2474 -393
rect 2512 -790 2796 -393
rect 2834 -790 2850 -393
rect 2458 -808 2850 -790
rect 3106 -393 3490 -382
rect 3106 -790 3118 -393
rect 3156 -790 3440 -393
rect 3478 -790 3490 -393
rect 3106 -804 3490 -790
rect 3750 -393 4134 -378
rect 3750 -790 3762 -393
rect 3800 -790 4084 -393
rect 4122 -790 4134 -393
rect 3750 -800 4134 -790
rect 4390 -393 4782 -374
rect 4390 -790 4406 -393
rect 4444 -790 4728 -393
rect 4766 -790 4782 -393
rect 4390 -808 4782 -790
rect 5034 -393 5426 -374
rect 5034 -790 5050 -393
rect 5088 -790 5372 -393
rect 5410 -790 5426 -393
rect 5034 -808 5426 -790
rect 5678 -393 6070 -374
rect 5678 -790 5694 -393
rect 5732 -790 6016 -393
rect 6054 -790 6070 -393
rect 5678 -808 6070 -790
rect 6322 -393 6714 -374
rect 6322 -790 6338 -393
rect 6376 -790 6660 -393
rect 6698 -790 6714 -393
rect 6322 -808 6714 -790
rect 6968 -393 7354 -380
rect 6968 -790 6982 -393
rect 7020 -790 7304 -393
rect 7342 -790 7354 -393
rect 6968 -804 7354 -790
rect 7610 -393 8002 -374
rect 7610 -790 7626 -393
rect 7664 -790 7948 -393
rect 7986 -790 8002 -393
rect 7610 -808 8002 -790
rect 204 -2200 596 -2182
rect 204 -2597 220 -2200
rect 258 -2597 542 -2200
rect 580 -2597 596 -2200
rect 204 -2616 596 -2597
rect 848 -2200 1240 -2182
rect 848 -2597 864 -2200
rect 902 -2597 1186 -2200
rect 1224 -2597 1240 -2200
rect 848 -2616 1240 -2597
rect 1492 -2200 1884 -2182
rect 1492 -2597 1508 -2200
rect 1546 -2597 1830 -2200
rect 1868 -2597 1884 -2200
rect 1492 -2616 1884 -2597
rect 2136 -2200 2528 -2182
rect 2136 -2597 2152 -2200
rect 2190 -2597 2474 -2200
rect 2512 -2597 2528 -2200
rect 2136 -2616 2528 -2597
rect 2780 -2200 3172 -2182
rect 2780 -2597 2796 -2200
rect 2834 -2597 3118 -2200
rect 3156 -2597 3172 -2200
rect 2780 -2616 3172 -2597
rect 3424 -2200 3816 -2182
rect 3424 -2597 3440 -2200
rect 3478 -2597 3762 -2200
rect 3800 -2597 3816 -2200
rect 3424 -2616 3816 -2597
rect 4068 -2200 4460 -2182
rect 4068 -2597 4084 -2200
rect 4122 -2597 4406 -2200
rect 4444 -2597 4460 -2200
rect 4068 -2616 4460 -2597
rect 4712 -2200 5104 -2182
rect 4712 -2597 4728 -2200
rect 4766 -2597 5050 -2200
rect 5088 -2597 5104 -2200
rect 4712 -2616 5104 -2597
rect 5356 -2200 5748 -2182
rect 5356 -2597 5372 -2200
rect 5410 -2597 5694 -2200
rect 5732 -2597 5748 -2200
rect 5356 -2616 5748 -2597
rect 6000 -2200 6392 -2182
rect 6000 -2597 6016 -2200
rect 6054 -2597 6338 -2200
rect 6376 -2597 6392 -2200
rect 6000 -2616 6392 -2597
rect 6644 -2200 7036 -2182
rect 6644 -2597 6660 -2200
rect 6698 -2597 6982 -2200
rect 7020 -2597 7036 -2200
rect 6644 -2616 7036 -2597
rect 7288 -2200 7680 -2182
rect 7288 -2597 7304 -2200
rect 7342 -2597 7626 -2200
rect 7664 -2597 7680 -2200
rect 7288 -2616 7680 -2597
rect 7936 -2200 8002 -2182
rect 7936 -2597 7948 -2200
rect 7986 -2597 8002 -2200
rect 7936 -2756 8002 -2597
rect 7192 -2788 8012 -2756
rect 7192 -2954 7240 -2788
rect 7964 -2954 8012 -2788
rect 7192 -2982 8012 -2954
<< via1 >>
rect 7252 2326 7974 2512
rect 7240 -2954 7964 -2788
<< metal2 >>
rect 7222 2512 8004 2532
rect 7222 2326 7252 2512
rect 7974 2326 8004 2512
rect 7222 2308 8004 2326
rect 7196 -2788 8006 -2760
rect 7196 -2954 7240 -2788
rect 7964 -2954 8006 -2788
rect 7196 -2992 8006 -2954
<< labels >>
rlabel metal1 8 -804 196 296 1 vcm
port 1 n
rlabel metal2 7212 -2982 7996 -2772 1 GND
port 2 n
rlabel metal2 7236 2316 7992 2520 1 VDD
port 3 n
rlabel psubdiffcont 432 -272 7976 -228 1 GND
port 2 n
<< end >>
