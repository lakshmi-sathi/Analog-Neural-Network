magic
tech sky130A
magscale 1 2
timestamp 1627668659
<< error_p >>
rect -845 373 -787 379
rect -653 373 -595 379
rect -461 373 -403 379
rect -269 373 -211 379
rect -77 373 -19 379
rect 115 373 173 379
rect 307 373 365 379
rect 499 373 557 379
rect 691 373 749 379
rect -845 339 -833 373
rect -653 339 -641 373
rect -461 339 -449 373
rect -269 339 -257 373
rect -77 339 -65 373
rect 115 339 127 373
rect 307 339 319 373
rect 499 339 511 373
rect 691 339 703 373
rect -845 333 -787 339
rect -653 333 -595 339
rect -461 333 -403 339
rect -269 333 -211 339
rect -77 333 -19 339
rect 115 333 173 339
rect 307 333 365 339
rect 499 333 557 339
rect 691 333 749 339
rect -749 71 -691 77
rect -557 71 -499 77
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect 595 71 653 77
rect 787 71 845 77
rect -749 37 -737 71
rect -557 37 -545 71
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect 595 37 607 71
rect 787 37 799 71
rect -749 31 -691 37
rect -557 31 -499 37
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect 595 31 653 37
rect 787 31 845 37
rect -749 -37 -691 -31
rect -557 -37 -499 -31
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect 595 -37 653 -31
rect 787 -37 845 -31
rect -749 -71 -737 -37
rect -557 -71 -545 -37
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect 595 -71 607 -37
rect 787 -71 799 -37
rect -749 -77 -691 -71
rect -557 -77 -499 -71
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect 595 -77 653 -71
rect 787 -77 845 -71
rect -845 -339 -787 -333
rect -653 -339 -595 -333
rect -461 -339 -403 -333
rect -269 -339 -211 -333
rect -77 -339 -19 -333
rect 115 -339 173 -333
rect 307 -339 365 -333
rect 499 -339 557 -333
rect 691 -339 749 -333
rect -845 -373 -833 -339
rect -653 -373 -641 -339
rect -461 -373 -449 -339
rect -269 -373 -257 -339
rect -77 -373 -65 -339
rect 115 -373 127 -339
rect 307 -373 319 -339
rect 499 -373 511 -339
rect 691 -373 703 -339
rect -845 -379 -787 -373
rect -653 -379 -595 -373
rect -461 -379 -403 -373
rect -269 -379 -211 -373
rect -77 -379 -19 -373
rect 115 -379 173 -373
rect 307 -379 365 -373
rect 499 -379 557 -373
rect 691 -379 749 -373
<< pwell >>
rect -1031 -511 1031 511
<< nmos >>
rect -831 109 -801 301
rect -735 109 -705 301
rect -639 109 -609 301
rect -543 109 -513 301
rect -447 109 -417 301
rect -351 109 -321 301
rect -255 109 -225 301
rect -159 109 -129 301
rect -63 109 -33 301
rect 33 109 63 301
rect 129 109 159 301
rect 225 109 255 301
rect 321 109 351 301
rect 417 109 447 301
rect 513 109 543 301
rect 609 109 639 301
rect 705 109 735 301
rect 801 109 831 301
rect -831 -301 -801 -109
rect -735 -301 -705 -109
rect -639 -301 -609 -109
rect -543 -301 -513 -109
rect -447 -301 -417 -109
rect -351 -301 -321 -109
rect -255 -301 -225 -109
rect -159 -301 -129 -109
rect -63 -301 -33 -109
rect 33 -301 63 -109
rect 129 -301 159 -109
rect 225 -301 255 -109
rect 321 -301 351 -109
rect 417 -301 447 -109
rect 513 -301 543 -109
rect 609 -301 639 -109
rect 705 -301 735 -109
rect 801 -301 831 -109
<< ndiff >>
rect -893 289 -831 301
rect -893 121 -881 289
rect -847 121 -831 289
rect -893 109 -831 121
rect -801 289 -735 301
rect -801 121 -785 289
rect -751 121 -735 289
rect -801 109 -735 121
rect -705 289 -639 301
rect -705 121 -689 289
rect -655 121 -639 289
rect -705 109 -639 121
rect -609 289 -543 301
rect -609 121 -593 289
rect -559 121 -543 289
rect -609 109 -543 121
rect -513 289 -447 301
rect -513 121 -497 289
rect -463 121 -447 289
rect -513 109 -447 121
rect -417 289 -351 301
rect -417 121 -401 289
rect -367 121 -351 289
rect -417 109 -351 121
rect -321 289 -255 301
rect -321 121 -305 289
rect -271 121 -255 289
rect -321 109 -255 121
rect -225 289 -159 301
rect -225 121 -209 289
rect -175 121 -159 289
rect -225 109 -159 121
rect -129 289 -63 301
rect -129 121 -113 289
rect -79 121 -63 289
rect -129 109 -63 121
rect -33 289 33 301
rect -33 121 -17 289
rect 17 121 33 289
rect -33 109 33 121
rect 63 289 129 301
rect 63 121 79 289
rect 113 121 129 289
rect 63 109 129 121
rect 159 289 225 301
rect 159 121 175 289
rect 209 121 225 289
rect 159 109 225 121
rect 255 289 321 301
rect 255 121 271 289
rect 305 121 321 289
rect 255 109 321 121
rect 351 289 417 301
rect 351 121 367 289
rect 401 121 417 289
rect 351 109 417 121
rect 447 289 513 301
rect 447 121 463 289
rect 497 121 513 289
rect 447 109 513 121
rect 543 289 609 301
rect 543 121 559 289
rect 593 121 609 289
rect 543 109 609 121
rect 639 289 705 301
rect 639 121 655 289
rect 689 121 705 289
rect 639 109 705 121
rect 735 289 801 301
rect 735 121 751 289
rect 785 121 801 289
rect 735 109 801 121
rect 831 289 893 301
rect 831 121 847 289
rect 881 121 893 289
rect 831 109 893 121
rect -893 -121 -831 -109
rect -893 -289 -881 -121
rect -847 -289 -831 -121
rect -893 -301 -831 -289
rect -801 -121 -735 -109
rect -801 -289 -785 -121
rect -751 -289 -735 -121
rect -801 -301 -735 -289
rect -705 -121 -639 -109
rect -705 -289 -689 -121
rect -655 -289 -639 -121
rect -705 -301 -639 -289
rect -609 -121 -543 -109
rect -609 -289 -593 -121
rect -559 -289 -543 -121
rect -609 -301 -543 -289
rect -513 -121 -447 -109
rect -513 -289 -497 -121
rect -463 -289 -447 -121
rect -513 -301 -447 -289
rect -417 -121 -351 -109
rect -417 -289 -401 -121
rect -367 -289 -351 -121
rect -417 -301 -351 -289
rect -321 -121 -255 -109
rect -321 -289 -305 -121
rect -271 -289 -255 -121
rect -321 -301 -255 -289
rect -225 -121 -159 -109
rect -225 -289 -209 -121
rect -175 -289 -159 -121
rect -225 -301 -159 -289
rect -129 -121 -63 -109
rect -129 -289 -113 -121
rect -79 -289 -63 -121
rect -129 -301 -63 -289
rect -33 -121 33 -109
rect -33 -289 -17 -121
rect 17 -289 33 -121
rect -33 -301 33 -289
rect 63 -121 129 -109
rect 63 -289 79 -121
rect 113 -289 129 -121
rect 63 -301 129 -289
rect 159 -121 225 -109
rect 159 -289 175 -121
rect 209 -289 225 -121
rect 159 -301 225 -289
rect 255 -121 321 -109
rect 255 -289 271 -121
rect 305 -289 321 -121
rect 255 -301 321 -289
rect 351 -121 417 -109
rect 351 -289 367 -121
rect 401 -289 417 -121
rect 351 -301 417 -289
rect 447 -121 513 -109
rect 447 -289 463 -121
rect 497 -289 513 -121
rect 447 -301 513 -289
rect 543 -121 609 -109
rect 543 -289 559 -121
rect 593 -289 609 -121
rect 543 -301 609 -289
rect 639 -121 705 -109
rect 639 -289 655 -121
rect 689 -289 705 -121
rect 639 -301 705 -289
rect 735 -121 801 -109
rect 735 -289 751 -121
rect 785 -289 801 -121
rect 735 -301 801 -289
rect 831 -121 893 -109
rect 831 -289 847 -121
rect 881 -289 893 -121
rect 831 -301 893 -289
<< ndiffc >>
rect -881 121 -847 289
rect -785 121 -751 289
rect -689 121 -655 289
rect -593 121 -559 289
rect -497 121 -463 289
rect -401 121 -367 289
rect -305 121 -271 289
rect -209 121 -175 289
rect -113 121 -79 289
rect -17 121 17 289
rect 79 121 113 289
rect 175 121 209 289
rect 271 121 305 289
rect 367 121 401 289
rect 463 121 497 289
rect 559 121 593 289
rect 655 121 689 289
rect 751 121 785 289
rect 847 121 881 289
rect -881 -289 -847 -121
rect -785 -289 -751 -121
rect -689 -289 -655 -121
rect -593 -289 -559 -121
rect -497 -289 -463 -121
rect -401 -289 -367 -121
rect -305 -289 -271 -121
rect -209 -289 -175 -121
rect -113 -289 -79 -121
rect -17 -289 17 -121
rect 79 -289 113 -121
rect 175 -289 209 -121
rect 271 -289 305 -121
rect 367 -289 401 -121
rect 463 -289 497 -121
rect 559 -289 593 -121
rect 655 -289 689 -121
rect 751 -289 785 -121
rect 847 -289 881 -121
<< psubdiff >>
rect -995 441 -899 475
rect 899 441 995 475
rect -995 379 -961 441
rect 961 379 995 441
rect -995 -441 -961 -379
rect 961 -441 995 -379
rect -995 -475 -899 -441
rect 899 -475 995 -441
<< psubdiffcont >>
rect -899 441 899 475
rect -995 -379 -961 379
rect 961 -379 995 379
rect -899 -475 899 -441
<< poly >>
rect -849 373 -783 389
rect -849 339 -833 373
rect -799 339 -783 373
rect -849 323 -783 339
rect -657 373 -591 389
rect -657 339 -641 373
rect -607 339 -591 373
rect -831 301 -801 323
rect -735 301 -705 327
rect -657 323 -591 339
rect -465 373 -399 389
rect -465 339 -449 373
rect -415 339 -399 373
rect -639 301 -609 323
rect -543 301 -513 327
rect -465 323 -399 339
rect -273 373 -207 389
rect -273 339 -257 373
rect -223 339 -207 373
rect -447 301 -417 323
rect -351 301 -321 327
rect -273 323 -207 339
rect -81 373 -15 389
rect -81 339 -65 373
rect -31 339 -15 373
rect -255 301 -225 323
rect -159 301 -129 327
rect -81 323 -15 339
rect 111 373 177 389
rect 111 339 127 373
rect 161 339 177 373
rect -63 301 -33 323
rect 33 301 63 327
rect 111 323 177 339
rect 303 373 369 389
rect 303 339 319 373
rect 353 339 369 373
rect 129 301 159 323
rect 225 301 255 327
rect 303 323 369 339
rect 495 373 561 389
rect 495 339 511 373
rect 545 339 561 373
rect 321 301 351 323
rect 417 301 447 327
rect 495 323 561 339
rect 687 373 753 389
rect 687 339 703 373
rect 737 339 753 373
rect 513 301 543 323
rect 609 301 639 327
rect 687 323 753 339
rect 705 301 735 323
rect 801 301 831 327
rect -831 83 -801 109
rect -735 87 -705 109
rect -753 71 -687 87
rect -639 83 -609 109
rect -543 87 -513 109
rect -753 37 -737 71
rect -703 37 -687 71
rect -753 21 -687 37
rect -561 71 -495 87
rect -447 83 -417 109
rect -351 87 -321 109
rect -561 37 -545 71
rect -511 37 -495 71
rect -561 21 -495 37
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 513 83 543 109
rect 609 87 639 109
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect 591 71 657 87
rect 705 83 735 109
rect 801 87 831 109
rect 591 37 607 71
rect 641 37 657 71
rect 591 21 657 37
rect 783 71 849 87
rect 783 37 799 71
rect 833 37 849 71
rect 783 21 849 37
rect -753 -37 -687 -21
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -831 -109 -801 -83
rect -753 -87 -687 -71
rect -561 -37 -495 -21
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -735 -109 -705 -87
rect -639 -109 -609 -83
rect -561 -87 -495 -71
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -543 -109 -513 -87
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 591 -37 657 -21
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 417 -109 447 -87
rect 513 -109 543 -83
rect 591 -87 657 -71
rect 783 -37 849 -21
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 609 -109 639 -87
rect 705 -109 735 -83
rect 783 -87 849 -71
rect 801 -109 831 -87
rect -831 -323 -801 -301
rect -849 -339 -783 -323
rect -735 -327 -705 -301
rect -639 -323 -609 -301
rect -849 -373 -833 -339
rect -799 -373 -783 -339
rect -849 -389 -783 -373
rect -657 -339 -591 -323
rect -543 -327 -513 -301
rect -447 -323 -417 -301
rect -657 -373 -641 -339
rect -607 -373 -591 -339
rect -657 -389 -591 -373
rect -465 -339 -399 -323
rect -351 -327 -321 -301
rect -255 -323 -225 -301
rect -465 -373 -449 -339
rect -415 -373 -399 -339
rect -465 -389 -399 -373
rect -273 -339 -207 -323
rect -159 -327 -129 -301
rect -63 -323 -33 -301
rect -273 -373 -257 -339
rect -223 -373 -207 -339
rect -273 -389 -207 -373
rect -81 -339 -15 -323
rect 33 -327 63 -301
rect 129 -323 159 -301
rect -81 -373 -65 -339
rect -31 -373 -15 -339
rect -81 -389 -15 -373
rect 111 -339 177 -323
rect 225 -327 255 -301
rect 321 -323 351 -301
rect 111 -373 127 -339
rect 161 -373 177 -339
rect 111 -389 177 -373
rect 303 -339 369 -323
rect 417 -327 447 -301
rect 513 -323 543 -301
rect 303 -373 319 -339
rect 353 -373 369 -339
rect 303 -389 369 -373
rect 495 -339 561 -323
rect 609 -327 639 -301
rect 705 -323 735 -301
rect 495 -373 511 -339
rect 545 -373 561 -339
rect 495 -389 561 -373
rect 687 -339 753 -323
rect 801 -327 831 -301
rect 687 -373 703 -339
rect 737 -373 753 -339
rect 687 -389 753 -373
<< polycont >>
rect -833 339 -799 373
rect -641 339 -607 373
rect -449 339 -415 373
rect -257 339 -223 373
rect -65 339 -31 373
rect 127 339 161 373
rect 319 339 353 373
rect 511 339 545 373
rect 703 339 737 373
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect -833 -373 -799 -339
rect -641 -373 -607 -339
rect -449 -373 -415 -339
rect -257 -373 -223 -339
rect -65 -373 -31 -339
rect 127 -373 161 -339
rect 319 -373 353 -339
rect 511 -373 545 -339
rect 703 -373 737 -339
<< locali >>
rect -995 441 -899 475
rect 899 441 995 475
rect -995 379 -961 441
rect 961 379 995 441
rect -849 339 -833 373
rect -799 339 -783 373
rect -657 339 -641 373
rect -607 339 -591 373
rect -465 339 -449 373
rect -415 339 -399 373
rect -273 339 -257 373
rect -223 339 -207 373
rect -81 339 -65 373
rect -31 339 -15 373
rect 111 339 127 373
rect 161 339 177 373
rect 303 339 319 373
rect 353 339 369 373
rect 495 339 511 373
rect 545 339 561 373
rect 687 339 703 373
rect 737 339 753 373
rect -881 289 -847 305
rect -881 105 -847 121
rect -785 289 -751 305
rect -785 105 -751 121
rect -689 289 -655 305
rect -689 105 -655 121
rect -593 289 -559 305
rect -593 105 -559 121
rect -497 289 -463 305
rect -497 105 -463 121
rect -401 289 -367 305
rect -401 105 -367 121
rect -305 289 -271 305
rect -305 105 -271 121
rect -209 289 -175 305
rect -209 105 -175 121
rect -113 289 -79 305
rect -113 105 -79 121
rect -17 289 17 305
rect -17 105 17 121
rect 79 289 113 305
rect 79 105 113 121
rect 175 289 209 305
rect 175 105 209 121
rect 271 289 305 305
rect 271 105 305 121
rect 367 289 401 305
rect 367 105 401 121
rect 463 289 497 305
rect 463 105 497 121
rect 559 289 593 305
rect 559 105 593 121
rect 655 289 689 305
rect 655 105 689 121
rect 751 289 785 305
rect 751 105 785 121
rect 847 289 881 305
rect 847 105 881 121
rect -753 37 -737 71
rect -703 37 -687 71
rect -561 37 -545 71
rect -511 37 -495 71
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect 591 37 607 71
rect 641 37 657 71
rect 783 37 799 71
rect 833 37 849 71
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 783 -71 799 -37
rect 833 -71 849 -37
rect -881 -121 -847 -105
rect -881 -305 -847 -289
rect -785 -121 -751 -105
rect -785 -305 -751 -289
rect -689 -121 -655 -105
rect -689 -305 -655 -289
rect -593 -121 -559 -105
rect -593 -305 -559 -289
rect -497 -121 -463 -105
rect -497 -305 -463 -289
rect -401 -121 -367 -105
rect -401 -305 -367 -289
rect -305 -121 -271 -105
rect -305 -305 -271 -289
rect -209 -121 -175 -105
rect -209 -305 -175 -289
rect -113 -121 -79 -105
rect -113 -305 -79 -289
rect -17 -121 17 -105
rect -17 -305 17 -289
rect 79 -121 113 -105
rect 79 -305 113 -289
rect 175 -121 209 -105
rect 175 -305 209 -289
rect 271 -121 305 -105
rect 271 -305 305 -289
rect 367 -121 401 -105
rect 367 -305 401 -289
rect 463 -121 497 -105
rect 463 -305 497 -289
rect 559 -121 593 -105
rect 559 -305 593 -289
rect 655 -121 689 -105
rect 655 -305 689 -289
rect 751 -121 785 -105
rect 751 -305 785 -289
rect 847 -121 881 -105
rect 847 -305 881 -289
rect -849 -373 -833 -339
rect -799 -373 -783 -339
rect -657 -373 -641 -339
rect -607 -373 -591 -339
rect -465 -373 -449 -339
rect -415 -373 -399 -339
rect -273 -373 -257 -339
rect -223 -373 -207 -339
rect -81 -373 -65 -339
rect -31 -373 -15 -339
rect 111 -373 127 -339
rect 161 -373 177 -339
rect 303 -373 319 -339
rect 353 -373 369 -339
rect 495 -373 511 -339
rect 545 -373 561 -339
rect 687 -373 703 -339
rect 737 -373 753 -339
rect -995 -441 -961 -379
rect 961 -441 995 -379
rect -995 -475 -899 -441
rect 899 -475 995 -441
<< viali >>
rect -833 339 -799 373
rect -641 339 -607 373
rect -449 339 -415 373
rect -257 339 -223 373
rect -65 339 -31 373
rect 127 339 161 373
rect 319 339 353 373
rect 511 339 545 373
rect 703 339 737 373
rect -881 121 -847 289
rect -785 121 -751 289
rect -689 121 -655 289
rect -593 121 -559 289
rect -497 121 -463 289
rect -401 121 -367 289
rect -305 121 -271 289
rect -209 121 -175 289
rect -113 121 -79 289
rect -17 121 17 289
rect 79 121 113 289
rect 175 121 209 289
rect 271 121 305 289
rect 367 121 401 289
rect 463 121 497 289
rect 559 121 593 289
rect 655 121 689 289
rect 751 121 785 289
rect 847 121 881 289
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect -881 -289 -847 -121
rect -785 -289 -751 -121
rect -689 -289 -655 -121
rect -593 -289 -559 -121
rect -497 -289 -463 -121
rect -401 -289 -367 -121
rect -305 -289 -271 -121
rect -209 -289 -175 -121
rect -113 -289 -79 -121
rect -17 -289 17 -121
rect 79 -289 113 -121
rect 175 -289 209 -121
rect 271 -289 305 -121
rect 367 -289 401 -121
rect 463 -289 497 -121
rect 559 -289 593 -121
rect 655 -289 689 -121
rect 751 -289 785 -121
rect 847 -289 881 -121
rect -833 -373 -799 -339
rect -641 -373 -607 -339
rect -449 -373 -415 -339
rect -257 -373 -223 -339
rect -65 -373 -31 -339
rect 127 -373 161 -339
rect 319 -373 353 -339
rect 511 -373 545 -339
rect 703 -373 737 -339
<< metal1 >>
rect -845 373 -787 379
rect -845 339 -833 373
rect -799 339 -787 373
rect -845 333 -787 339
rect -653 373 -595 379
rect -653 339 -641 373
rect -607 339 -595 373
rect -653 333 -595 339
rect -461 373 -403 379
rect -461 339 -449 373
rect -415 339 -403 373
rect -461 333 -403 339
rect -269 373 -211 379
rect -269 339 -257 373
rect -223 339 -211 373
rect -269 333 -211 339
rect -77 373 -19 379
rect -77 339 -65 373
rect -31 339 -19 373
rect -77 333 -19 339
rect 115 373 173 379
rect 115 339 127 373
rect 161 339 173 373
rect 115 333 173 339
rect 307 373 365 379
rect 307 339 319 373
rect 353 339 365 373
rect 307 333 365 339
rect 499 373 557 379
rect 499 339 511 373
rect 545 339 557 373
rect 499 333 557 339
rect 691 373 749 379
rect 691 339 703 373
rect 737 339 749 373
rect 691 333 749 339
rect -887 289 -841 301
rect -887 121 -881 289
rect -847 121 -841 289
rect -887 109 -841 121
rect -791 289 -745 301
rect -791 121 -785 289
rect -751 121 -745 289
rect -791 109 -745 121
rect -695 289 -649 301
rect -695 121 -689 289
rect -655 121 -649 289
rect -695 109 -649 121
rect -599 289 -553 301
rect -599 121 -593 289
rect -559 121 -553 289
rect -599 109 -553 121
rect -503 289 -457 301
rect -503 121 -497 289
rect -463 121 -457 289
rect -503 109 -457 121
rect -407 289 -361 301
rect -407 121 -401 289
rect -367 121 -361 289
rect -407 109 -361 121
rect -311 289 -265 301
rect -311 121 -305 289
rect -271 121 -265 289
rect -311 109 -265 121
rect -215 289 -169 301
rect -215 121 -209 289
rect -175 121 -169 289
rect -215 109 -169 121
rect -119 289 -73 301
rect -119 121 -113 289
rect -79 121 -73 289
rect -119 109 -73 121
rect -23 289 23 301
rect -23 121 -17 289
rect 17 121 23 289
rect -23 109 23 121
rect 73 289 119 301
rect 73 121 79 289
rect 113 121 119 289
rect 73 109 119 121
rect 169 289 215 301
rect 169 121 175 289
rect 209 121 215 289
rect 169 109 215 121
rect 265 289 311 301
rect 265 121 271 289
rect 305 121 311 289
rect 265 109 311 121
rect 361 289 407 301
rect 361 121 367 289
rect 401 121 407 289
rect 361 109 407 121
rect 457 289 503 301
rect 457 121 463 289
rect 497 121 503 289
rect 457 109 503 121
rect 553 289 599 301
rect 553 121 559 289
rect 593 121 599 289
rect 553 109 599 121
rect 649 289 695 301
rect 649 121 655 289
rect 689 121 695 289
rect 649 109 695 121
rect 745 289 791 301
rect 745 121 751 289
rect 785 121 791 289
rect 745 109 791 121
rect 841 289 887 301
rect 841 121 847 289
rect 881 121 887 289
rect 841 109 887 121
rect -749 71 -691 77
rect -749 37 -737 71
rect -703 37 -691 71
rect -749 31 -691 37
rect -557 71 -499 77
rect -557 37 -545 71
rect -511 37 -499 71
rect -557 31 -499 37
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect 595 71 653 77
rect 595 37 607 71
rect 641 37 653 71
rect 595 31 653 37
rect 787 71 845 77
rect 787 37 799 71
rect 833 37 845 71
rect 787 31 845 37
rect -749 -37 -691 -31
rect -749 -71 -737 -37
rect -703 -71 -691 -37
rect -749 -77 -691 -71
rect -557 -37 -499 -31
rect -557 -71 -545 -37
rect -511 -71 -499 -37
rect -557 -77 -499 -71
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect 595 -37 653 -31
rect 595 -71 607 -37
rect 641 -71 653 -37
rect 595 -77 653 -71
rect 787 -37 845 -31
rect 787 -71 799 -37
rect 833 -71 845 -37
rect 787 -77 845 -71
rect -887 -121 -841 -109
rect -887 -289 -881 -121
rect -847 -289 -841 -121
rect -887 -301 -841 -289
rect -791 -121 -745 -109
rect -791 -289 -785 -121
rect -751 -289 -745 -121
rect -791 -301 -745 -289
rect -695 -121 -649 -109
rect -695 -289 -689 -121
rect -655 -289 -649 -121
rect -695 -301 -649 -289
rect -599 -121 -553 -109
rect -599 -289 -593 -121
rect -559 -289 -553 -121
rect -599 -301 -553 -289
rect -503 -121 -457 -109
rect -503 -289 -497 -121
rect -463 -289 -457 -121
rect -503 -301 -457 -289
rect -407 -121 -361 -109
rect -407 -289 -401 -121
rect -367 -289 -361 -121
rect -407 -301 -361 -289
rect -311 -121 -265 -109
rect -311 -289 -305 -121
rect -271 -289 -265 -121
rect -311 -301 -265 -289
rect -215 -121 -169 -109
rect -215 -289 -209 -121
rect -175 -289 -169 -121
rect -215 -301 -169 -289
rect -119 -121 -73 -109
rect -119 -289 -113 -121
rect -79 -289 -73 -121
rect -119 -301 -73 -289
rect -23 -121 23 -109
rect -23 -289 -17 -121
rect 17 -289 23 -121
rect -23 -301 23 -289
rect 73 -121 119 -109
rect 73 -289 79 -121
rect 113 -289 119 -121
rect 73 -301 119 -289
rect 169 -121 215 -109
rect 169 -289 175 -121
rect 209 -289 215 -121
rect 169 -301 215 -289
rect 265 -121 311 -109
rect 265 -289 271 -121
rect 305 -289 311 -121
rect 265 -301 311 -289
rect 361 -121 407 -109
rect 361 -289 367 -121
rect 401 -289 407 -121
rect 361 -301 407 -289
rect 457 -121 503 -109
rect 457 -289 463 -121
rect 497 -289 503 -121
rect 457 -301 503 -289
rect 553 -121 599 -109
rect 553 -289 559 -121
rect 593 -289 599 -121
rect 553 -301 599 -289
rect 649 -121 695 -109
rect 649 -289 655 -121
rect 689 -289 695 -121
rect 649 -301 695 -289
rect 745 -121 791 -109
rect 745 -289 751 -121
rect 785 -289 791 -121
rect 745 -301 791 -289
rect 841 -121 887 -109
rect 841 -289 847 -121
rect 881 -289 887 -121
rect 841 -301 887 -289
rect -845 -339 -787 -333
rect -845 -373 -833 -339
rect -799 -373 -787 -339
rect -845 -379 -787 -373
rect -653 -339 -595 -333
rect -653 -373 -641 -339
rect -607 -373 -595 -339
rect -653 -379 -595 -373
rect -461 -339 -403 -333
rect -461 -373 -449 -339
rect -415 -373 -403 -339
rect -461 -379 -403 -373
rect -269 -339 -211 -333
rect -269 -373 -257 -339
rect -223 -373 -211 -339
rect -269 -379 -211 -373
rect -77 -339 -19 -333
rect -77 -373 -65 -339
rect -31 -373 -19 -339
rect -77 -379 -19 -373
rect 115 -339 173 -333
rect 115 -373 127 -339
rect 161 -373 173 -339
rect 115 -379 173 -373
rect 307 -339 365 -333
rect 307 -373 319 -339
rect 353 -373 365 -339
rect 307 -379 365 -373
rect 499 -339 557 -333
rect 499 -373 511 -339
rect 545 -373 557 -339
rect 499 -379 557 -373
rect 691 -339 749 -333
rect 691 -373 703 -339
rect 737 -373 749 -339
rect 691 -379 749 -373
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -978 -458 978 458
string parameters w 0.96 l 0.150 m 2 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
